
module FDE_Rex_Runner ( clk, rstn, start_i, db_o, dori_o, cs_o, en_o, rw_o, 
        rst_o, state );
  output [7:0] db_o;
  output [3:0] cs_o;
  output [2:0] state;
  input clk, rstn, start_i;
  output dori_o, en_o, rw_o, rst_o;
  wire   \driver/N96 , \driver/N47 , \driver/N46 , \driver/N45 , \driver/N44 ,
         \driver/*Logic0* , \decider/N96 , \decider/N95 , \decider/N94 ,
         \decider/N93 , \decider/N92 , \decider/N91 , \decider/N90 ,
         \decider/N89 , \decider/N88 , \decider/N85 , \decider/N84 ,
         \decider/N83 , \decider/N82 , \decider/N81 , \decider/N80 ,
         \decider/N79 , \decider/N78 , \decider/N77 , \decider/N64 ,
         \decider/N63 , \decider/N62 , \decider/N61 , \decider/N60 ,
         \decider/N58 , \decider/N57 , \decider/N55 , \decider/N38 ,
         \decider/posx_m_obstacle_right[15] , \decider/posy_m_rex_top[1] ,
         \decider/posy_m_rex_top[2] , \decider/posy_m_rex_top[3] ,
         \decider/posy_m_rex_top[4] , \decider/posy_m_rex_top[5] , n376, n377,
         n378, n379, n380, n381, n403, n404, n405, n406, n407, n408, n409,
         n410, n411, n412, n413, n414, n415, n416, n417, n418, n419, n420,
         n421, n422, n423, n424, \r50/carry[9] , \r50/carry[8] ,
         \r50/carry[7] , \r50/carry[6] , \r50/carry[5] , \r50/carry[4] ,
         \r50/carry[3] , \r50/carry[2] , \r50/carry[1] ,
         \add_2_root_decider/add_109_3_cf/carry[2] ,
         \add_2_root_decider/add_109_3_cf/carry[3] ,
         \add_2_root_decider/add_109_3_cf/carry[4] ,
         \add_2_root_decider/add_109_3_cf/carry[6] ,
         \add_2_root_decider/add_109_3_cf/carry[7] , \r61/PROD1[4] ,
         \r61/SUMB[1][2] , \r61/SUMB[1][3] , \r61/SUMB[2][2] ,
         \r61/SUMB[2][3] , \r61/SUMB[3][2] , \r61/SUMB[3][3] ,
         \r61/SUMB[4][2] , \r61/SUMB[4][3] , \r61/SUMB[5][2] ,
         \r61/SUMB[5][3] , \r61/SUMB[6][2] , \r61/SUMB[6][3] ,
         \r61/SUMB[7][2] , \r61/CARRYB[2][2] , \r61/CARRYB[2][3] ,
         \r61/CARRYB[3][0] , \r61/CARRYB[3][2] , \r61/CARRYB[3][3] ,
         \r61/CARRYB[4][0] , \r61/CARRYB[4][2] , \r61/CARRYB[4][3] ,
         \r61/CARRYB[5][2] , \r61/CARRYB[6][2] , \r61/ab[0][2] ,
         \r61/ab[1][0] , \r61/ab[1][2] , \r61/ab[2][0] , \r61/ab[2][2] ,
         \r61/ab[3][0] , \r61/ab[3][2] , \r61/ab[4][0] , \r61/ab[4][2] ,
         \r61/ab[7][2] , \sub_1_root_decider/sub_49/carry[2] ,
         \sub_1_root_decider/sub_49/carry[3] ,
         \sub_1_root_decider/sub_49/carry[5] ,
         \sub_1_root_decider/sub_49/carry[6] , \decider/sub_45/carry[2] ,
         \decider/sub_45/carry[3] , \decider/sub_45/carry[4] ,
         \decider/sub_45/carry[5] , \decider/sub_75/carry[6] ,
         \decider/sub_75/carry[5] , \sub_0_root_decider/sub_73/carry[15] ,
         \r180/carry[8] , \r180/carry[7] , n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n499,
         n500, n501, n502, n503, n504, n505, n506, n507, n508, n509, n510,
         n511, n512, n513, n514, n515, n516, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551, n552, n553, n554,
         n555, n556, n557, n558, n559, n560, n561, n562, n563, n564, n565,
         n566, n567, n568, n569, n570, n571, n572, n573, n574, n575, n576,
         n577, n578, n579, n580, n581, n582, n583, n584, n585, n586, n587,
         n588, n589, n590, n591, n592, n593, n594, n595, n596, n597, n598,
         n599, n600, n601, n602, n603, n604, n605, n606, n607, n608, n609,
         n610, n611, n612, n613, n614, n615, n616, n617, n618, n619, n620,
         n621, n622, n623, n624, n625, n626, n627, n628, n629, n630, n631,
         n632, n633, n634, n635, n636, n637, n638, n639, n640, n641, n642,
         n643, n644, n645, n646, n647, n648, n649, n650, n651, n652, n653,
         n654, n655, n656, n657, n658, n659, n660, n661, n662, n663, n664,
         n665, n666, n667, n668, n669, n670, n671, n672, n673, n674, n675,
         n676, n677, n678, n679, n680, n681, n682, n683, n684, n685, n686,
         n687, n688, n689, n690, n691, n692, n693, n694;
  wire   [10:0] addrD;
  wire   [15:0] addrT;
  wire   [1:0] \driver/start_history ;
  wire   [5:0] \decider/posy_m_obstacle_top ;
  wire   [15:0] \decider/obstacle_right ;
  wire   [7:3] \decider/posx_m_rex_left ;
  assign rw_o = \driver/*Logic0* ;

  DFFHQ \driver/en_o_reg  ( .D(\driver/N96 ), .CK(clk), .Q(en_o) );
  DFFHQ \driver/rst_o_reg  ( .D(n661), .CK(clk), .Q(rst_o) );
  EDFFHQ \driver/start_history_reg[0]  ( .D(start_i), .E(rstn), .CK(clk), .Q(
        \driver/start_history [0]) );
  EDFFHQ \driver/start_history_reg[1]  ( .D(\driver/start_history [0]), .E(
        rstn), .CK(clk), .Q(\driver/start_history [1]) );
  DFFHQ \driver/x_reg[2]  ( .D(n415), .CK(clk), .Q(addrD[8]) );
  DFFHQ \driver/x_reg[0]  ( .D(n417), .CK(clk), .Q(addrD[6]) );
  DFFHQ \driver/x_reg[1]  ( .D(n416), .CK(clk), .Q(addrD[7]) );
  DFFHQ \driver/x_reg[3]  ( .D(n414), .CK(clk), .Q(addrD[9]) );
  DFFHQ \driver/x_reg[4]  ( .D(n418), .CK(clk), .Q(addrD[10]) );
  DFFHQ \driver/state_reg[0]  ( .D(n412), .CK(clk), .Q(state[0]) );
  DFFHQ \driver/state_reg[1]  ( .D(n411), .CK(clk), .Q(state[1]) );
  DFFHQ \driver/state_reg[2]  ( .D(n413), .CK(clk), .Q(state[2]) );
  DFFHQ \driver/y_reg[5]  ( .D(n424), .CK(clk), .Q(addrD[5]) );
  DFFHQ \driver/y_reg[0]  ( .D(n423), .CK(clk), .Q(addrD[0]) );
  DFFHQ \driver/y_reg[1]  ( .D(n422), .CK(clk), .Q(addrD[1]) );
  DFFHQ \driver/y_reg[2]  ( .D(n421), .CK(clk), .Q(addrD[2]) );
  DFFHQ \driver/y_reg[3]  ( .D(n420), .CK(clk), .Q(addrD[3]) );
  DFFHQ \driver/y_reg[4]  ( .D(n419), .CK(clk), .Q(addrD[4]) );
  DFFHQ \driver/dori_o_reg  ( .D(n410), .CK(clk), .Q(dori_o) );
  DFFRHQ \decider/addrT_reg[0]  ( .D(n663), .CK(clk), .RN(rstn), .Q(addrT[0])
         );
  DFFRHQ \decider/addrT_reg[1]  ( .D(n664), .CK(clk), .RN(rstn), .Q(addrT[1])
         );
  DFFRHQ \decider/addrT_reg[2]  ( .D(n665), .CK(clk), .RN(rstn), .Q(addrT[2])
         );
  DFFRHQ \decider/addrT_reg[3]  ( .D(n666), .CK(clk), .RN(rstn), .Q(addrT[3])
         );
  DFFRHQ \decider/addrT_reg[4]  ( .D(n667), .CK(clk), .RN(rstn), .Q(addrT[4])
         );
  DFFRHQ \decider/addrT_reg[5]  ( .D(n668), .CK(clk), .RN(rstn), .Q(addrT[5])
         );
  DFFRHQ \decider/addrT_reg[6]  ( .D(n669), .CK(clk), .RN(rstn), .Q(addrT[6])
         );
  DFFRHQ \decider/addrT_reg[7]  ( .D(n670), .CK(clk), .RN(rstn), .Q(addrT[7])
         );
  DFFRHQ \decider/addrT_reg[8]  ( .D(n671), .CK(clk), .RN(rstn), .Q(addrT[8])
         );
  DFFRHQ \decider/addrT_reg[9]  ( .D(n672), .CK(clk), .RN(rstn), .Q(addrT[9])
         );
  DFFHQ \driver/db_o_reg[6]  ( .D(n403), .CK(clk), .Q(db_o[6]) );
  DFFHQ \driver/db_o_reg[5]  ( .D(n404), .CK(clk), .Q(db_o[5]) );
  DFFHQ \driver/db_o_reg[4]  ( .D(n405), .CK(clk), .Q(db_o[4]) );
  DFFHQ \driver/db_o_reg[3]  ( .D(n406), .CK(clk), .Q(db_o[3]) );
  DFFHQ \driver/db_o_reg[2]  ( .D(n407), .CK(clk), .Q(db_o[2]) );
  DFFHQ \driver/db_o_reg[1]  ( .D(n408), .CK(clk), .Q(db_o[1]) );
  DFFHQ \driver/db_o_reg[0]  ( .D(n409), .CK(clk), .Q(db_o[0]) );
  DFFHQ \driver/db_o_reg[7]  ( .D(n662), .CK(clk), .Q(db_o[7]) );
  ADDF \r50/U2_1  ( .A(n685), .B(n380), .CI(\r50/carry[1] ), .CO(
        \r50/carry[2] ), .S(\decider/N88 ) );
  ADDF \r50/U2_2  ( .A(n683), .B(n379), .CI(\r50/carry[2] ), .CO(
        \r50/carry[3] ), .S(\decider/N89 ) );
  ADDF \r50/U2_3  ( .A(n681), .B(n378), .CI(\r50/carry[3] ), .CO(
        \r50/carry[4] ), .S(\decider/N90 ) );
  ADDF \r50/U2_4  ( .A(n679), .B(n377), .CI(\r50/carry[4] ), .CO(
        \r50/carry[5] ), .S(\decider/N91 ) );
  ADDF \r50/U2_5  ( .A(n677), .B(n376), .CI(\r50/carry[5] ), .CO(
        \r50/carry[6] ), .S(\decider/N92 ) );
  ADDF \r50/U2_6  ( .A(n676), .B(n688), .CI(\r50/carry[6] ), .CO(
        \r50/carry[7] ), .S(\decider/N93 ) );
  ADDF \r50/U2_7  ( .A(n675), .B(n688), .CI(\r50/carry[7] ), .CO(
        \r50/carry[8] ), .S(\decider/N94 ) );
  ADDF \r50/U2_8  ( .A(n674), .B(n688), .CI(\r50/carry[8] ), .CO(
        \r50/carry[9] ), .S(\decider/N95 ) );
  ADDF \r50/U2_9  ( .A(n673), .B(n688), .CI(\r50/carry[9] ), .S(\decider/N96 )
         );
  ADDF \r61/S3_2_3  ( .A(n684), .B(n443), .CI(n687), .CO(\r61/CARRYB[2][3] ), 
        .S(\r61/SUMB[2][3] ) );
  ADDF \r61/S2_2_2  ( .A(\r61/ab[2][2] ), .B(n442), .CI(\r61/SUMB[1][3] ), 
        .CO(\r61/CARRYB[2][2] ), .S(\r61/SUMB[2][2] ) );
  ADDF \r61/S3_3_3  ( .A(n682), .B(\r61/CARRYB[2][3] ), .CI(n684), .CO(
        \r61/CARRYB[3][3] ), .S(\r61/SUMB[3][3] ) );
  ADDF \r61/S2_3_2  ( .A(\r61/ab[3][2] ), .B(\r61/CARRYB[2][2] ), .CI(
        \r61/SUMB[2][3] ), .CO(\r61/CARRYB[3][2] ), .S(\r61/SUMB[3][2] ) );
  ADDF \r61/S1_3_0  ( .A(\r61/ab[3][0] ), .B(n441), .CI(\r61/SUMB[1][2] ), 
        .CO(\r61/CARRYB[3][0] ), .S(\decider/N58 ) );
  ADDF \r61/S3_4_3  ( .A(n680), .B(\r61/CARRYB[3][3] ), .CI(n682), .CO(
        \r61/CARRYB[4][3] ), .S(\r61/SUMB[4][3] ) );
  ADDF \r61/S2_4_2  ( .A(\r61/ab[4][2] ), .B(\r61/CARRYB[3][2] ), .CI(
        \r61/SUMB[3][3] ), .CO(\r61/CARRYB[4][2] ), .S(\r61/SUMB[4][2] ) );
  ADDF \r61/S1_4_0  ( .A(\r61/ab[4][0] ), .B(\r61/CARRYB[3][0] ), .CI(
        \r61/SUMB[2][2] ), .CO(\r61/CARRYB[4][0] ), .S(\r61/PROD1[4] ) );
  ADDF \r61/S3_5_3  ( .A(\r61/ab[7][2] ), .B(\r61/CARRYB[4][3] ), .CI(n680), 
        .CO(\r61/SUMB[6][3] ), .S(\r61/SUMB[5][3] ) );
  ADDF \r61/S2_5_2  ( .A(\r61/ab[7][2] ), .B(\r61/CARRYB[4][2] ), .CI(
        \r61/SUMB[4][3] ), .CO(\r61/CARRYB[5][2] ), .S(\r61/SUMB[5][2] ) );
  ADDF \r61/S2_6_2  ( .A(\r61/ab[7][2] ), .B(\r61/CARRYB[5][2] ), .CI(
        \r61/SUMB[5][3] ), .CO(\r61/CARRYB[6][2] ), .S(\r61/SUMB[6][2] ) );
  ADDF \r61/S2_7_2  ( .A(\r61/ab[7][2] ), .B(\r61/CARRYB[6][2] ), .CI(
        \r61/SUMB[6][3] ), .S(\r61/SUMB[7][2] ) );
  AND2 U325 ( .A(addrD[7]), .B(addrD[6]), .Y(n428) );
  AND2 U326 ( .A(addrD[8]), .B(n428), .Y(n429) );
  AND2 U327 ( .A(\add_2_root_decider/add_109_3_cf/carry[4] ), .B(
        \r61/PROD1[4] ), .Y(n430) );
  AND2 U328 ( .A(n693), .B(\sub_1_root_decider/sub_49/carry[3] ), .Y(n431) );
  OR2 U329 ( .A(n486), .B(addrT[6]), .Y(n432) );
  AND2 U330 ( .A(\add_2_root_decider/add_109_3_cf/carry[7] ), .B(\decider/N62 ), .Y(n433) );
  AND2 U331 ( .A(n693), .B(n692), .Y(n434) );
  AND2 U332 ( .A(\r61/CARRYB[4][0] ), .B(\r61/SUMB[3][2] ), .Y(n435) );
  AND2 U333 ( .A(n435), .B(\r61/SUMB[4][2] ), .Y(n436) );
  AND2 U334 ( .A(n436), .B(\r61/SUMB[5][2] ), .Y(n437) );
  AND2 U335 ( .A(addrD[9]), .B(n429), .Y(n438) );
  AND2 U336 ( .A(n433), .B(\decider/N63 ), .Y(n439) );
  AND2 U337 ( .A(n437), .B(\r61/SUMB[6][2] ), .Y(n440) );
  AND2 U338 ( .A(\r61/ab[2][0] ), .B(\r61/ab[0][2] ), .Y(n441) );
  AND2 U339 ( .A(n460), .B(\r61/ab[1][2] ), .Y(n442) );
  AND2 U340 ( .A(n460), .B(n687), .Y(n443) );
  INV U341 ( .A(n589), .Y(n444) );
  BUF U342 ( .I(n488), .O(n445) );
  INV U343 ( .A(n529), .Y(n446) );
  BUF U344 ( .I(n469), .O(n447) );
  BUF U345 ( .I(n469), .O(n448) );
  LOGIC_0 U346 ( .LOGIC_0_PIN(\driver/*Logic0* ) );
  NAND2 U347 ( .A(n449), .B(n450), .Y(\r50/carry[1] ) );
  XNOR2 U348 ( .A(n381), .B(n686), .Y(\decider/N38 ) );
  INV U349 ( .A(n381), .Y(n449) );
  INV U350 ( .A(n686), .Y(n450) );
  NAND2 U351 ( .A(n451), .B(n452), .Y(
        \add_2_root_decider/add_109_3_cf/carry[2] ) );
  XNOR2 U352 ( .A(\r61/ab[1][0] ), .B(\decider/N55 ), .Y(\decider/N85 ) );
  INV U353 ( .A(\r61/ab[1][0] ), .Y(n451) );
  INV U354 ( .A(\decider/N55 ), .Y(n452) );
  NAND2 U355 ( .A(n453), .B(n462), .Y(
        \add_2_root_decider/add_109_3_cf/carry[4] ) );
  XNOR2 U356 ( .A(\decider/N58 ), .B(
        \add_2_root_decider/add_109_3_cf/carry[3] ), .Y(\decider/N83 ) );
  INV U357 ( .A(\decider/N58 ), .Y(n453) );
  NAND2 U358 ( .A(n454), .B(n463), .Y(
        \add_2_root_decider/add_109_3_cf/carry[7] ) );
  XNOR2 U359 ( .A(\decider/N61 ), .B(
        \add_2_root_decider/add_109_3_cf/carry[6] ), .Y(\decider/N80 ) );
  INV U360 ( .A(\decider/N61 ), .Y(n454) );
  NAND2 U361 ( .A(addrD[1]), .B(addrD[0]), .Y(
        \sub_1_root_decider/sub_49/carry[2] ) );
  XNOR2 U362 ( .A(n691), .B(n690), .Y(\decider/posy_m_rex_top[1] ) );
  NAND2 U363 ( .A(addrD[2]), .B(n455), .Y(\sub_1_root_decider/sub_49/carry[3] ) );
  XNOR2 U364 ( .A(n692), .B(\sub_1_root_decider/sub_49/carry[2] ), .Y(
        \decider/posy_m_rex_top[2] ) );
  INV U365 ( .A(\sub_1_root_decider/sub_49/carry[2] ), .Y(n455) );
  NAND2 U366 ( .A(addrD[5]), .B(n464), .Y(\sub_1_root_decider/sub_49/carry[6] ) );
  XNOR2 U367 ( .A(n689), .B(\sub_1_root_decider/sub_49/carry[5] ), .Y(
        \decider/posy_m_rex_top[5] ) );
  NAND2 U368 ( .A(n509), .B(n456), .Y(\decider/sub_45/carry[5] ) );
  XNOR2 U369 ( .A(addrD[10]), .B(\decider/sub_45/carry[4] ), .Y(
        \decider/posx_m_rex_left [7]) );
  INV U370 ( .A(\decider/sub_45/carry[4] ), .Y(n456) );
  NAND2 U371 ( .A(n457), .B(n458), .Y(\decider/sub_45/carry[4] ) );
  XNOR2 U372 ( .A(addrD[9]), .B(\decider/sub_45/carry[3] ), .Y(
        \decider/posx_m_rex_left [6]) );
  INV U373 ( .A(addrD[9]), .Y(n457) );
  INV U374 ( .A(\decider/sub_45/carry[3] ), .Y(n458) );
  NAND2 U375 ( .A(n513), .B(n459), .Y(\decider/sub_45/carry[3] ) );
  XNOR2 U376 ( .A(addrD[8]), .B(\decider/sub_45/carry[2] ), .Y(
        \decider/posx_m_rex_left [5]) );
  INV U377 ( .A(\decider/sub_45/carry[2] ), .Y(n459) );
  NAND2 U378 ( .A(n512), .B(n460), .Y(\decider/sub_45/carry[2] ) );
  XNOR2 U379 ( .A(addrD[7]), .B(addrD[6]), .Y(\decider/posx_m_rex_left [4]) );
  INV U380 ( .A(addrD[6]), .Y(n460) );
  NAND2 U381 ( .A(addrD[5]), .B(n465), .Y(\decider/sub_75/carry[6] ) );
  XNOR2 U382 ( .A(n689), .B(\decider/sub_75/carry[5] ), .Y(
        \decider/posy_m_obstacle_top [5]) );
  XNOR2 U383 ( .A(n678), .B(\sub_0_root_decider/sub_73/carry[15] ), .Y(
        \decider/posx_m_obstacle_right[15] ) );
  NAND2 U384 ( .A(n457), .B(n466), .Y(\r180/carry[7] ) );
  XNOR2 U385 ( .A(addrD[9]), .B(n429), .Y(\decider/obstacle_right [6]) );
  NAND2 U386 ( .A(n509), .B(n461), .Y(\r180/carry[8] ) );
  XNOR2 U387 ( .A(addrD[10]), .B(\r180/carry[7] ), .Y(
        \decider/obstacle_right [7]) );
  INV U388 ( .A(\r180/carry[7] ), .Y(n461) );
  XOR2 U389 ( .A(addrD[7]), .B(addrD[6]), .Y(\driver/N44 ) );
  XOR2 U390 ( .A(addrD[8]), .B(n428), .Y(\driver/N45 ) );
  XOR2 U391 ( .A(addrD[9]), .B(n429), .Y(\driver/N46 ) );
  XOR2 U392 ( .A(addrD[10]), .B(n438), .Y(\driver/N47 ) );
  XOR2 U393 ( .A(\decider/N57 ), .B(\add_2_root_decider/add_109_3_cf/carry[2] ), .Y(\decider/N84 ) );
  NAND2 U394 ( .A(\add_2_root_decider/add_109_3_cf/carry[2] ), .B(
        \decider/N57 ), .Y(n462) );
  INV U395 ( .A(n462), .Y(\add_2_root_decider/add_109_3_cf/carry[3] ) );
  XOR2 U396 ( .A(\r61/PROD1[4] ), .B(
        \add_2_root_decider/add_109_3_cf/carry[4] ), .Y(\decider/N82 ) );
  XOR2 U397 ( .A(\decider/N60 ), .B(n430), .Y(\decider/N81 ) );
  NAND2 U398 ( .A(n430), .B(\decider/N60 ), .Y(n463) );
  INV U399 ( .A(n463), .Y(\add_2_root_decider/add_109_3_cf/carry[6] ) );
  XOR2 U400 ( .A(\decider/N62 ), .B(\add_2_root_decider/add_109_3_cf/carry[7] ), .Y(\decider/N79 ) );
  XOR2 U401 ( .A(\decider/N63 ), .B(n433), .Y(\decider/N78 ) );
  XOR2 U402 ( .A(\decider/N64 ), .B(n439), .Y(\decider/N77 ) );
  XOR2 U403 ( .A(\r61/ab[1][2] ), .B(n460), .Y(\r61/SUMB[1][2] ) );
  XOR2 U404 ( .A(n687), .B(n460), .Y(\r61/SUMB[1][3] ) );
  XOR2 U405 ( .A(n693), .B(\sub_1_root_decider/sub_49/carry[3] ), .Y(
        \decider/posy_m_rex_top[3] ) );
  XOR2 U406 ( .A(n694), .B(n431), .Y(\decider/posy_m_rex_top[4] ) );
  NAND2 U407 ( .A(n694), .B(n431), .Y(n464) );
  INV U408 ( .A(n464), .Y(\sub_1_root_decider/sub_49/carry[5] ) );
  XOR2 U409 ( .A(n693), .B(n692), .Y(\decider/posy_m_obstacle_top [3]) );
  XOR2 U410 ( .A(n694), .B(n434), .Y(\decider/posy_m_obstacle_top [4]) );
  NAND2 U411 ( .A(n694), .B(n434), .Y(n465) );
  INV U412 ( .A(n465), .Y(\decider/sub_75/carry[5] ) );
  XOR2 U413 ( .A(addrD[7]), .B(addrD[6]), .Y(\decider/obstacle_right [4]) );
  XOR2 U414 ( .A(addrD[8]), .B(n428), .Y(\decider/obstacle_right [5]) );
  NAND2 U415 ( .A(addrD[8]), .B(n428), .Y(n466) );
  XOR2 U416 ( .A(\r61/ab[2][0] ), .B(\r61/ab[0][2] ), .Y(\decider/N57 ) );
  XOR2 U417 ( .A(\r61/CARRYB[4][0] ), .B(\r61/SUMB[3][2] ), .Y(\decider/N60 )
         );
  XOR2 U418 ( .A(n435), .B(\r61/SUMB[4][2] ), .Y(\decider/N61 ) );
  XOR2 U419 ( .A(n436), .B(\r61/SUMB[5][2] ), .Y(\decider/N62 ) );
  XOR2 U420 ( .A(n437), .B(\r61/SUMB[6][2] ), .Y(\decider/N63 ) );
  XOR2 U421 ( .A(n440), .B(\r61/SUMB[7][2] ), .Y(\decider/N64 ) );
  INV U422 ( .A(n467), .Y(\sub_0_root_decider/sub_73/carry[15] ) );
  NOR4BB U423 ( .AN(n468), .BN(\r180/carry[8] ), .C(
        \decider/obstacle_right [5]), .D(\decider/obstacle_right [4]), .Y(n467) );
  NOR2 U424 ( .A(\decider/obstacle_right [7]), .B(\decider/obstacle_right [6]), 
        .Y(n468) );
  NOR2B U425 ( .AN(n680), .B(n448), .Y(\r61/ab[4][2] ) );
  NOR2B U426 ( .AN(n680), .B(n470), .Y(\r61/ab[4][0] ) );
  NOR2B U427 ( .AN(n682), .B(n447), .Y(\r61/ab[3][2] ) );
  NOR2B U428 ( .AN(n682), .B(n470), .Y(\r61/ab[3][0] ) );
  NOR2B U429 ( .AN(n684), .B(n448), .Y(\r61/ab[2][2] ) );
  NOR2B U430 ( .AN(n684), .B(n470), .Y(\r61/ab[2][0] ) );
  NOR2B U431 ( .AN(n687), .B(n447), .Y(\r61/ab[1][2] ) );
  NOR2B U432 ( .AN(n460), .B(n448), .Y(\r61/ab[0][2] ) );
  INV U433 ( .A(n471), .Y(n662) );
  AOI221 U434 ( .A0(db_o[7]), .A1(n472), .B0(n473), .B1(n474), .C0(n475), .Y(
        n471) );
  OAI211 U435 ( .A0(n476), .A1(n477), .B0(n478), .C0(n479), .Y(n474) );
  AOI221 U436 ( .A0(addrT[3]), .A1(n480), .B0(n481), .B1(n482), .C0(n483), .Y(
        n479) );
  NOR2B U437 ( .AN(n484), .B(addrT[1]), .Y(n481) );
  OAI21 U438 ( .A0(n485), .A1(n486), .B0(n487), .Y(n480) );
  MX2 U439 ( .A(\decider/N38 ), .B(addrT[0]), .S0(n445), .Y(n663) );
  MX2 U440 ( .A(\decider/N88 ), .B(addrT[1]), .S0(n445), .Y(n664) );
  MX2 U441 ( .A(\decider/N89 ), .B(addrT[2]), .S0(n445), .Y(n665) );
  MX2 U442 ( .A(\decider/N90 ), .B(addrT[3]), .S0(n445), .Y(n666) );
  MX2 U443 ( .A(\decider/N91 ), .B(addrT[4]), .S0(n445), .Y(n667) );
  MX2 U444 ( .A(\decider/N92 ), .B(addrT[5]), .S0(n445), .Y(n668) );
  MX2 U445 ( .A(\decider/N93 ), .B(addrT[6]), .S0(n445), .Y(n669) );
  MX2 U446 ( .A(\decider/N94 ), .B(addrT[7]), .S0(n445), .Y(n670) );
  MX2 U447 ( .A(\decider/N95 ), .B(addrT[8]), .S0(n445), .Y(n671) );
  MX2 U448 ( .A(\decider/N96 ), .B(addrT[9]), .S0(n445), .Y(n672) );
  AOI31 U449 ( .A0(\decider/posx_m_obstacle_right[15] ), .A1(n489), .A2(
        \r180/carry[8] ), .B0(n447), .Y(n488) );
  INV U450 ( .A(\decider/sub_75/carry[6] ), .Y(n489) );
  MX2 U451 ( .A(\decider/N77 ), .B(\decider/N64 ), .S0(n448), .Y(n673) );
  MX2 U452 ( .A(\decider/N78 ), .B(\decider/N63 ), .S0(n447), .Y(n674) );
  MX2 U453 ( .A(\decider/N79 ), .B(\decider/N62 ), .S0(n448), .Y(n675) );
  MX2 U454 ( .A(\decider/N80 ), .B(\decider/N61 ), .S0(n447), .Y(n676) );
  MX2 U455 ( .A(\decider/N81 ), .B(\decider/N60 ), .S0(n448), .Y(n677) );
  MX2 U456 ( .A(\decider/N82 ), .B(\r61/PROD1[4] ), .S0(n447), .Y(n679) );
  MX2 U457 ( .A(\decider/obstacle_right [7]), .B(\decider/posx_m_rex_left [7]), 
        .S0(n448), .Y(n680) );
  MX2 U458 ( .A(\decider/N83 ), .B(\decider/N58 ), .S0(n447), .Y(n681) );
  MX2 U459 ( .A(\decider/obstacle_right [6]), .B(\decider/posx_m_rex_left [6]), 
        .S0(n448), .Y(n682) );
  MX2 U460 ( .A(\decider/N84 ), .B(\decider/N57 ), .S0(n447), .Y(n683) );
  MX2 U461 ( .A(\decider/obstacle_right [5]), .B(\decider/posx_m_rex_left [5]), 
        .S0(n448), .Y(n684) );
  OAI2BB1 U462 ( .A0N(\decider/N85 ), .A1N(n470), .B0(n451), .Y(n685) );
  NOR2B U463 ( .AN(n687), .B(n470), .Y(\r61/ab[1][0] ) );
  INV U464 ( .A(n448), .Y(n470) );
  NAND2 U465 ( .A(addrD[6]), .B(n447), .Y(n686) );
  MX2 U466 ( .A(\decider/obstacle_right [4]), .B(\decider/posx_m_rex_left [4]), 
        .S0(n447), .Y(n687) );
  NOR2B U467 ( .AN(\decider/sub_75/carry[6] ), .B(n448), .Y(n688) );
  MX2 U468 ( .A(n490), .B(n491), .S0(addrD[5]), .Y(n424) );
  OAI21 U469 ( .A0(addrD[4]), .A1(n492), .B0(n493), .Y(n491) );
  NOR2B U470 ( .AN(n494), .B(n495), .Y(n490) );
  MX2 U471 ( .A(n494), .B(n496), .S0(addrD[0]), .Y(n423) );
  MX2 U472 ( .A(n497), .B(n498), .S0(addrD[1]), .Y(n422) );
  INV U473 ( .A(n499), .Y(n498) );
  NOR2B U474 ( .AN(addrD[0]), .B(n492), .Y(n497) );
  MX2 U475 ( .A(n500), .B(n501), .S0(addrD[2]), .Y(n421) );
  OAI21 U476 ( .A0(addrD[1]), .A1(n492), .B0(n499), .Y(n501) );
  AOI2BB1 U477 ( .A0N(addrD[0]), .A1N(n492), .B0(n496), .Y(n499) );
  NOR3B U478 ( .AN(addrD[1]), .B(n492), .C(n690), .Y(n500) );
  MX2 U479 ( .A(n502), .B(n503), .S0(addrD[3]), .Y(n420) );
  NOR2B U480 ( .AN(n504), .B(n492), .Y(n502) );
  MX2 U481 ( .A(n505), .B(n506), .S0(addrD[4]), .Y(n419) );
  INV U482 ( .A(n493), .Y(n506) );
  AOI2BB1 U483 ( .A0N(addrD[3]), .A1N(n492), .B0(n503), .Y(n493) );
  OAI21 U484 ( .A0(n504), .A1(n492), .B0(n507), .Y(n503) );
  INV U485 ( .A(n496), .Y(n507) );
  NOR3B U486 ( .AN(n504), .B(n492), .C(n693), .Y(n505) );
  OAI2BB2 U487 ( .B0(n508), .B1(n509), .A0N(\driver/N47 ), .A1N(n510), .Y(n418) );
  MX2 U488 ( .A(n510), .B(n511), .S0(addrD[6]), .Y(n417) );
  OAI2BB2 U489 ( .B0(n508), .B1(n512), .A0N(\driver/N44 ), .A1N(n510), .Y(n416) );
  OAI2BB2 U490 ( .B0(n508), .B1(n513), .A0N(\driver/N45 ), .A1N(n510), .Y(n415) );
  OAI2BB2 U491 ( .B0(n508), .B1(n457), .A0N(\driver/N46 ), .A1N(n510), .Y(n414) );
  NOR2B U492 ( .AN(n514), .B(n511), .Y(n510) );
  INV U493 ( .A(n508), .Y(n511) );
  OAI2BB1 U494 ( .A0N(state[2]), .A1N(n515), .B0(n516), .Y(n413) );
  NAND2 U495 ( .A(n517), .B(n516), .Y(n412) );
  MX2 U496 ( .A(n518), .B(n519), .S0(n515), .Y(n517) );
  AOI31 U497 ( .A0(cs_o[3]), .A1(addrD[8]), .A2(n520), .B0(n521), .Y(n518) );
  NOR3B U498 ( .AN(addrD[7]), .B(n460), .C(n522), .Y(n520) );
  INV U499 ( .A(n523), .Y(n411) );
  NOR3B U500 ( .AN(n516), .B(n524), .C(n525), .Y(n523) );
  MX2 U501 ( .A(n526), .B(state[1]), .S0(n446), .Y(n525) );
  OAI31 U502 ( .A0(n527), .A1(n661), .A2(n528), .B0(n529), .Y(n516) );
  INV U503 ( .A(n515), .Y(n529) );
  AOI211 U504 ( .A0(en_o), .A1(n527), .B0(n530), .C0(n508), .Y(n515) );
  OAI31 U505 ( .A0(n531), .A1(n689), .A2(n495), .B0(n532), .Y(n508) );
  INV U506 ( .A(n533), .Y(n495) );
  NOR3B U507 ( .AN(n504), .B(n693), .C(n694), .Y(n533) );
  NOR3B U508 ( .AN(addrD[1]), .B(n690), .C(n692), .Y(n504) );
  INV U509 ( .A(addrD[2]), .Y(n692) );
  NOR2B U510 ( .AN(state[2]), .B(n534), .Y(n527) );
  OAI2BB1 U511 ( .A0N(n535), .A1N(dori_o), .B0(n492), .Y(n410) );
  INV U512 ( .A(n494), .Y(n492) );
  NOR2B U513 ( .AN(n514), .B(n496), .Y(n494) );
  NOR2B U514 ( .AN(rstn), .B(n522), .Y(n514) );
  NOR2B U515 ( .AN(n496), .B(n530), .Y(n535) );
  INV U516 ( .A(n536), .Y(n530) );
  NOR2B U517 ( .AN(n532), .B(n537), .Y(n496) );
  AOI31 U518 ( .A0(n538), .A1(n524), .A2(\driver/start_history [1]), .B0(n661), 
        .Y(n532) );
  INV U519 ( .A(rstn), .Y(n661) );
  NOR2B U520 ( .AN(en_o), .B(start_i), .Y(n538) );
  INV U521 ( .A(n539), .Y(n409) );
  AOI221 U522 ( .A0(n528), .A1(n540), .B0(db_o[0]), .B1(n472), .C0(n541), .Y(
        n539) );
  OAI222 U523 ( .A0(n542), .A1(n543), .B0(n460), .B1(n544), .C0(n690), .C1(
        n545), .Y(n541) );
  INV U524 ( .A(addrD[0]), .Y(n690) );
  NOR3B U525 ( .AN(n546), .B(n547), .C(n548), .Y(n542) );
  MX2 U526 ( .A(n549), .B(n550), .S0(n444), .Y(n548) );
  NOR2B U527 ( .AN(n551), .B(n477), .Y(n550) );
  NOR3B U528 ( .AN(n552), .B(addrT[4]), .C(n485), .Y(n549) );
  AOI32 U529 ( .A0(n553), .A1(n554), .A2(n555), .B0(n556), .B1(n557), .Y(n546)
         );
  OAI22 U530 ( .A0(n558), .A1(n559), .B0(n560), .B1(n561), .Y(n557) );
  NOR2B U531 ( .AN(n562), .B(addrT[0]), .Y(n560) );
  AOI21 U532 ( .A0(addrT[3]), .A1(addrT[1]), .B0(addrT[6]), .Y(n558) );
  INV U533 ( .A(n563), .Y(n408) );
  AOI221 U534 ( .A0(n564), .A1(addrD[1]), .B0(db_o[1]), .B1(n472), .C0(n565), 
        .Y(n563) );
  OAI221 U535 ( .A0(n512), .A1(n544), .B0(n566), .B1(n543), .C0(n567), .Y(n565) );
  NOR4 U536 ( .A(n568), .B(n569), .C(n547), .D(n570), .Y(n566) );
  OAI2BB2 U537 ( .B0(n571), .B1(n572), .A0N(n573), .A1N(n556), .Y(n570) );
  OAI2BB1 U538 ( .A0N(addrT[4]), .A1N(n574), .B0(n561), .Y(n573) );
  OAI21 U539 ( .A0(addrT[0]), .A1(n575), .B0(n576), .Y(n574) );
  INV U540 ( .A(addrT[6]), .Y(n576) );
  AOI21 U541 ( .A0(n562), .A1(n577), .B0(n578), .Y(n571) );
  OAI21 U542 ( .A0(addrT[3]), .A1(n579), .B0(n580), .Y(n547) );
  OAI33 U543 ( .A0(n581), .A1(n432), .A2(n582), .B0(n579), .B1(addrT[2]), .B2(
        n583), .Y(n569) );
  OAI31 U544 ( .A0(n487), .A1(addrT[3]), .A2(n485), .B0(n584), .Y(n568) );
  INV U545 ( .A(addrD[7]), .Y(n512) );
  INV U546 ( .A(n585), .Y(n407) );
  AOI221 U547 ( .A0(n564), .A1(addrD[2]), .B0(db_o[2]), .B1(n472), .C0(n586), 
        .Y(n585) );
  OAI221 U548 ( .A0(n513), .A1(n544), .B0(n587), .B1(n543), .C0(n567), .Y(n586) );
  INV U549 ( .A(n588), .Y(n587) );
  OAI221 U550 ( .A0(n589), .A1(n590), .B0(n591), .B1(addrT[2]), .C0(n592), .Y(
        n588) );
  AOI211 U551 ( .A0(n589), .A1(n593), .B0(n483), .C0(n555), .Y(n591) );
  NOR2B U552 ( .AN(n594), .B(n582), .Y(n483) );
  AOI32 U553 ( .A0(n562), .A1(n559), .A2(n595), .B0(addrT[1]), .B1(n593), .Y(
        n590) );
  INV U554 ( .A(addrD[8]), .Y(n513) );
  OAI221 U555 ( .A0(n596), .A1(n543), .B0(n693), .B1(n545), .C0(n597), .Y(n406) );
  AOI21 U556 ( .A0(db_o[3]), .A1(n472), .B0(n598), .Y(n597) );
  INV U557 ( .A(addrD[3]), .Y(n693) );
  NOR4BB U558 ( .AN(n599), .BN(n579), .C(n600), .D(n601), .Y(n596) );
  OAI211 U559 ( .A0(n602), .A1(n582), .B0(n592), .C0(n603), .Y(n601) );
  AOI32 U560 ( .A0(n575), .A1(n554), .A2(n604), .B0(n605), .B1(n606), .Y(n603)
         );
  OAI2BB2 U561 ( .B0(n432), .B1(n581), .A0N(n607), .A1N(n593), .Y(n605) );
  INV U562 ( .A(n608), .Y(n592) );
  OAI221 U563 ( .A0(n609), .A1(n580), .B0(addrT[3]), .B1(n610), .C0(n611), .Y(
        n608) );
  NOR2 U564 ( .A(n612), .B(n613), .Y(n611) );
  INV U565 ( .A(n604), .Y(n610) );
  NAND3 U566 ( .A(addrT[3]), .B(n556), .C(addrT[2]), .Y(n580) );
  AOI2BB2 U567 ( .B0(addrT[4]), .B1(n477), .A0N(n553), .A1N(addrT[6]), .Y(n609) );
  AOI33 U568 ( .A0(n577), .A1(n552), .A2(n485), .B0(addrT[3]), .B1(n583), .B2(
        n593), .Y(n599) );
  NOR2B U569 ( .AN(addrT[2]), .B(n477), .Y(n485) );
  OAI221 U570 ( .A0(n614), .A1(n543), .B0(n694), .B1(n545), .C0(n615), .Y(n405) );
  AOI21 U571 ( .A0(db_o[4]), .A1(n472), .B0(n598), .Y(n615) );
  INV U572 ( .A(addrD[4]), .Y(n694) );
  NOR4B U573 ( .AN(n616), .B(n612), .C(n600), .D(n617), .Y(n614) );
  OAI221 U574 ( .A0(n618), .A1(n579), .B0(n619), .B1(n581), .C0(n620), .Y(n617) );
  NOR2B U575 ( .AN(n621), .B(n622), .Y(n619) );
  XOR2 U576 ( .A(addrT[3]), .B(n575), .Y(n618) );
  OAI211 U577 ( .A0(n623), .A1(n624), .B0(n625), .C0(n484), .Y(n616) );
  NOR3B U578 ( .AN(n477), .B(n554), .C(n559), .Y(n623) );
  INV U579 ( .A(n583), .Y(n477) );
  OAI221 U580 ( .A0(n626), .A1(n543), .B0(n689), .B1(n545), .C0(n627), .Y(n404) );
  AOI21 U581 ( .A0(db_o[5]), .A1(n472), .B0(n598), .Y(n627) );
  NAND2 U582 ( .A(n544), .B(n567), .Y(n598) );
  OR2 U583 ( .A(n628), .B(n629), .Y(n567) );
  AOI31 U584 ( .A0(\driver/start_history [1]), .A1(n630), .A2(n524), .B0(n528), 
        .Y(n628) );
  INV U585 ( .A(start_i), .Y(n630) );
  INV U586 ( .A(n475), .Y(n544) );
  NOR2B U587 ( .AN(n631), .B(n629), .Y(n475) );
  INV U588 ( .A(addrD[5]), .Y(n689) );
  NOR3 U589 ( .A(n632), .B(n633), .C(n634), .Y(n626) );
  MX2 U590 ( .A(n600), .B(n635), .S0(addrT[0]), .Y(n634) );
  NOR3B U591 ( .AN(addrT[2]), .B(n476), .C(addrT[1]), .Y(n635) );
  INV U592 ( .A(n594), .Y(n476) );
  AND3 U593 ( .A(n607), .B(n575), .C(n593), .Y(n600) );
  NOR2B U594 ( .AN(n551), .B(n559), .Y(n593) );
  OAI2BB2 U595 ( .B0(n621), .B1(n581), .A0N(addrT[3]), .A1N(n636), .Y(n632) );
  OAI221 U596 ( .A0(n637), .A1(n487), .B0(n582), .B1(n579), .C0(n638), .Y(n636) );
  AOI31 U597 ( .A0(n583), .A1(n559), .A2(n551), .B0(n639), .Y(n638) );
  INV U598 ( .A(n640), .Y(n639) );
  AOI31 U599 ( .A0(n594), .A1(n606), .A2(addrT[1]), .B0(n622), .Y(n640) );
  NOR3 U600 ( .A(addrT[1]), .B(n572), .C(n559), .Y(n622) );
  NOR2 U601 ( .A(n486), .B(n559), .Y(n594) );
  INV U602 ( .A(n555), .Y(n579) );
  NOR2B U603 ( .AN(n554), .B(n582), .Y(n637) );
  INV U604 ( .A(n553), .Y(n582) );
  AOI2BB1 U605 ( .A0N(addrT[0]), .A1N(n432), .B0(n555), .Y(n621) );
  NOR2B U606 ( .AN(n559), .B(n432), .Y(n555) );
  OAI221 U607 ( .A0(n641), .A1(n543), .B0(n642), .B1(n643), .C0(n545), .Y(n403) );
  INV U608 ( .A(n564), .Y(n545) );
  NOR2B U609 ( .AN(n521), .B(n629), .Y(n564) );
  INV U610 ( .A(n540), .Y(n629) );
  INV U611 ( .A(db_o[6]), .Y(n643) );
  INV U612 ( .A(n473), .Y(n543) );
  NOR4 U613 ( .A(addrT[9]), .B(addrT[8]), .C(\r61/ab[7][2] ), .D(n644), .Y(
        n473) );
  OAI211 U614 ( .A0(n447), .A1(n645), .B0(n526), .C0(n540), .Y(n644) );
  NOR2B U615 ( .AN(rstn), .B(n472), .Y(n540) );
  INV U616 ( .A(n642), .Y(n472) );
  OAI211 U617 ( .A0(n646), .A1(\driver/N96 ), .B0(n536), .C0(n531), .Y(n642)
         );
  INV U618 ( .A(n537), .Y(n531) );
  NOR2B U619 ( .AN(en_o), .B(n522), .Y(n537) );
  INV U620 ( .A(n526), .Y(n522) );
  OAI31 U621 ( .A0(n631), .A1(n528), .A2(n521), .B0(en_o), .Y(n536) );
  NOR3B U622 ( .AN(state[1]), .B(state[0]), .C(state[2]), .Y(n521) );
  NOR2B U623 ( .AN(n534), .B(state[2]), .Y(n528) );
  NOR3 U624 ( .A(n519), .B(state[1]), .C(state[2]), .Y(n631) );
  NOR2B U625 ( .AN(rstn), .B(n524), .Y(n646) );
  AND2 U626 ( .A(n534), .B(state[2]), .Y(n524) );
  NOR2B U627 ( .AN(state[1]), .B(n519), .Y(n534) );
  NOR3B U628 ( .AN(n519), .B(state[1]), .C(state[2]), .Y(n526) );
  INV U629 ( .A(state[0]), .Y(n519) );
  NOR2B U630 ( .AN(\decider/posx_m_obstacle_right[15] ), .B(
        \decider/sub_75/carry[6] ), .Y(n645) );
  AOI2BB1 U631 ( .A0N(n647), .A1N(n589), .B0(n633), .Y(n641) );
  OAI211 U632 ( .A0(n648), .A1(n572), .B0(n478), .C0(n620), .Y(n633) );
  AOI31 U633 ( .A0(n577), .A1(addrT[2]), .A2(n551), .B0(n613), .Y(n620) );
  NOR2B U634 ( .AN(n583), .B(n602), .Y(n613) );
  NOR2B U635 ( .AN(n559), .B(n589), .Y(n577) );
  NOR3B U636 ( .AN(n584), .B(n604), .C(n649), .Y(n478) );
  NOR4BB U637 ( .AN(addrT[7]), .BN(n482), .C(n583), .D(addrT[6]), .Y(n649) );
  NOR3B U638 ( .AN(n607), .B(addrT[5]), .C(addrT[4]), .Y(n482) );
  NOR2B U639 ( .AN(n554), .B(addrT[3]), .Y(n607) );
  NOR2B U640 ( .AN(addrT[4]), .B(n487), .Y(n604) );
  INV U641 ( .A(n595), .Y(n487) );
  INV U642 ( .A(n612), .Y(n584) );
  NOR2B U643 ( .AN(addrT[2]), .B(n602), .Y(n612) );
  INV U644 ( .A(n650), .Y(n602) );
  NOR2B U645 ( .AN(n589), .B(n432), .Y(n650) );
  INV U646 ( .A(n552), .Y(n486) );
  AOI2BB1 U647 ( .A0N(n554), .A1N(n561), .B0(n624), .Y(n648) );
  OAI2BB2 U648 ( .B0(n559), .B1(n581), .A0N(n583), .A1N(n578), .Y(n624) );
  NOR2B U649 ( .AN(addrT[0]), .B(n575), .Y(n583) );
  INV U650 ( .A(addrT[1]), .Y(n575) );
  NAND2B U651 ( .AN(addrT[2]), .B(addrT[3]), .Y(n581) );
  INV U652 ( .A(addrT[4]), .Y(n559) );
  INV U653 ( .A(n578), .Y(n561) );
  NOR2B U654 ( .AN(addrT[4]), .B(addrT[3]), .Y(n578) );
  INV U655 ( .A(addrT[3]), .Y(n589) );
  AOI211 U656 ( .A0(n552), .A1(n651), .B0(n652), .C0(n595), .Y(n647) );
  NOR2B U657 ( .AN(addrT[5]), .B(n572), .Y(n595) );
  MX2 U658 ( .A(n653), .B(n654), .S0(addrT[4]), .Y(n652) );
  NOR2B U659 ( .AN(n553), .B(n572), .Y(n654) );
  INV U660 ( .A(n484), .Y(n572) );
  NOR2B U661 ( .AN(addrT[6]), .B(addrT[7]), .Y(n484) );
  NOR2B U662 ( .AN(n551), .B(n553), .Y(n653) );
  NOR2B U663 ( .AN(n606), .B(addrT[1]), .Y(n553) );
  INV U664 ( .A(addrT[0]), .Y(n606) );
  NOR2B U665 ( .AN(n556), .B(addrT[6]), .Y(n551) );
  NOR2B U666 ( .AN(n625), .B(addrT[7]), .Y(n556) );
  INV U667 ( .A(addrT[5]), .Y(n625) );
  OAI21 U668 ( .A0(n562), .A1(addrT[4]), .B0(n655), .Y(n651) );
  MX2 U669 ( .A(addrT[2]), .B(addrT[1]), .S0(addrT[0]), .Y(n655) );
  NOR2B U670 ( .AN(addrT[1]), .B(n554), .Y(n562) );
  INV U671 ( .A(addrT[2]), .Y(n554) );
  NOR2B U672 ( .AN(addrT[5]), .B(addrT[7]), .Y(n552) );
  XOR2 U673 ( .A(addrD[0]), .B(n448), .Y(n381) );
  INV U674 ( .A(n656), .Y(n380) );
  MX2 U675 ( .A(n691), .B(\decider/posy_m_rex_top[1] ), .S0(n447), .Y(n656) );
  INV U676 ( .A(addrD[1]), .Y(n691) );
  INV U677 ( .A(n657), .Y(n379) );
  MX2 U678 ( .A(addrD[2]), .B(\decider/posy_m_rex_top[2] ), .S0(n448), .Y(n657) );
  INV U679 ( .A(n658), .Y(n378) );
  MX2 U680 ( .A(\decider/posy_m_obstacle_top [3]), .B(
        \decider/posy_m_rex_top[3] ), .S0(n447), .Y(n658) );
  INV U681 ( .A(n659), .Y(n377) );
  MX2 U682 ( .A(\decider/posy_m_obstacle_top [4]), .B(
        \decider/posy_m_rex_top[4] ), .S0(n448), .Y(n659) );
  INV U683 ( .A(n660), .Y(n376) );
  MX2 U684 ( .A(\decider/posy_m_obstacle_top [5]), .B(
        \decider/posy_m_rex_top[5] ), .S0(n447), .Y(n660) );
  NOR2B U685 ( .AN(rstn), .B(en_o), .Y(\driver/N96 ) );
  NOR2B U686 ( .AN(n448), .B(addrD[6]), .Y(\decider/N55 ) );
  NOR2B U687 ( .AN(addrD[10]), .B(n457), .Y(cs_o[3]) );
  NOR2B U688 ( .AN(addrD[10]), .B(addrD[9]), .Y(cs_o[2]) );
  NOR2B U689 ( .AN(n509), .B(n457), .Y(cs_o[1]) );
  NOR2B U690 ( .AN(n678), .B(n447), .Y(\r61/ab[7][2] ) );
  NOR4BB U691 ( .AN(\decider/sub_45/carry[5] ), .BN(cs_o[0]), .C(addrD[8]), 
        .D(\sub_1_root_decider/sub_49/carry[6] ), .Y(n469) );
  NOR2B U692 ( .AN(n509), .B(addrD[9]), .Y(cs_o[0]) );
  INV U693 ( .A(addrD[10]), .Y(n509) );
  INV U694 ( .A(\r180/carry[8] ), .Y(n678) );
endmodule

