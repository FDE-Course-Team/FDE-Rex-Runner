module Decider(
    
);



endmodule