
module FDE_Rex_Runner ( clk, rstn, start_i, db_o, dori_o, cs_o, en_o, rw_o, 
        rst_o, state );
  output [7:0] db_o;
  output [3:0] cs_o;
  output [2:0] state;
  input clk, rstn, start_i;
  output dori_o, en_o, rw_o, rst_o;
  wire   \driver/N96 , \driver/N47 , \driver/N46 , \driver/N45 , \driver/N44 ,
         \driver/*Logic0* , \decider/N96 , \decider/N95 , \decider/N94 ,
         \decider/N93 , \decider/N92 , \decider/N91 , \decider/N90 ,
         \decider/N89 , \decider/N88 , \decider/N85 , \decider/N84 ,
         \decider/N83 , \decider/N82 , \decider/N81 , \decider/N80 ,
         \decider/N79 , \decider/N78 , \decider/N77 , \decider/N64 ,
         \decider/N63 , \decider/N62 , \decider/N61 , \decider/N60 ,
         \decider/N58 , \decider/N57 , \decider/N56 , \decider/N55 ,
         \decider/N38 , \decider/posx_m_obstacle_right[15] ,
         \decider/posy_m_rex_top[1] , \decider/posy_m_rex_top[2] ,
         \decider/posy_m_rex_top[3] , \decider/posy_m_rex_top[4] ,
         \decider/posy_m_rex_top[5] , \U3/U1/Z_1 , \U3/U1/Z_2 , \U3/U1/Z_3 ,
         \U3/U1/Z_4 , \U3/U1/Z_8 , \U3/U3/Z_0 , \U3/U3/Z_1 , \U3/U3/Z_2 ,
         \U3/U3/Z_3 , \U3/U3/Z_4 , \U3/U3/Z_5 , \U3/U3/Z_6 , \U3/U3/Z_7 ,
         \U3/U3/Z_8 , \U3/U3/Z_9 , n352, n353, n354, n355, n356, n357, n358,
         n359, n360, n361, n362, n363, n364, n365, n366, n367, n368, n369,
         n370, n371, n372, n373, \r50/carry[9] , \r50/carry[8] ,
         \r50/carry[7] , \r50/carry[6] , \r50/carry[5] , \r50/carry[4] ,
         \r50/carry[3] , \r50/carry[2] , \r50/carry[1] ,
         \add_2_root_decider/add_109_3_cf/carry[2] ,
         \add_2_root_decider/add_109_3_cf/carry[3] ,
         \add_2_root_decider/add_109_3_cf/carry[6] ,
         \add_2_root_decider/add_109_3_cf/carry[7] , \r61/PROD1[4] ,
         \r61/SUMB[1][1] , \r61/SUMB[2][1] , \r61/SUMB[2][2] ,
         \r61/SUMB[3][1] , \r61/SUMB[3][2] , \r61/SUMB[4][1] ,
         \r61/SUMB[4][2] , \r61/SUMB[5][1] , \r61/SUMB[5][2] ,
         \r61/SUMB[6][1] , \r61/SUMB[6][2] , \r61/SUMB[7][1] ,
         \r61/SUMB[7][2] , \r61/SUMB[8][1] , \r61/CARRYB[2][0] ,
         \r61/CARRYB[2][1] , \r61/CARRYB[3][0] , \r61/CARRYB[3][1] ,
         \r61/CARRYB[3][2] , \r61/CARRYB[4][0] , \r61/CARRYB[4][1] ,
         \r61/CARRYB[4][2] , \r61/CARRYB[5][1] , \r61/CARRYB[5][2] ,
         \r61/CARRYB[6][1] , \r61/CARRYB[7][1] , \r61/ab[1][0] ,
         \r61/ab[2][0] , \r61/ab[3][0] , \r61/ab[4][0] ,
         \sub_1_root_decider/sub_49/carry[3] ,
         \sub_1_root_decider/sub_49/carry[4] ,
         \sub_1_root_decider/sub_49/carry[5] ,
         \sub_1_root_decider/sub_49/carry[6] , \decider/sub_45/carry[2] ,
         \decider/sub_45/carry[3] , \decider/sub_45/carry[4] ,
         \decider/sub_45/carry[5] , \decider/sub_75/carry[6] ,
         \decider/sub_75/carry[4] , \sub_0_root_decider/sub_73/carry[15] ,
         \r180/carry[8] , \r180/carry[7] , n377, n378, n379, n380, n381, n382,
         n383, n384, n385, n386, n387, n388, n389, n390, n391, n392, n393,
         n394, n395, n396, n397, n398, n399, n400, n401, n402, n403, n404,
         n405, n406, n407, n408, n409, n410, n411, n412, n413, n414, n415,
         n416, n417, n418, n419, n420, n421, n422, n423, n424, n425, n426,
         n427, n428, n429, n430, n431, n432, n433, n434, n435, n436, n437,
         n438, n439, n440, n441, n442, n443, n444, n445, n446, n447, n448,
         n449, n450, n451, n452, n453, n454, n455, n456, n457, n458, n459,
         n460, n461, n462, n463, n464, n465, n466, n467, n468, n469, n470,
         n471, n472, n473, n474, n475, n476, n477, n478, n479, n480, n481,
         n482, n483, n484, n485, n486, n487, n488, n489, n490, n491, n492,
         n493, n494, n495, n496, n497, n498, n499, n500, n501, n502, n503,
         n504, n505, n506, n507, n508, n509, n510, n511, n512, n513, n514,
         n515, n516, n517, n518, n519, n520, n521, n522, n523, n524, n525,
         n526, n527, n528, n529, n530, n531, n532, n533, n534, n535, n536,
         n537, n538, n539, n540, n541, n542, n543, n544, n545, n546, n547,
         n548, n549, n550, n551, n552, n553, n554, n555, n556, n557, n558,
         n559, n560, n561, n562, n563, n564, n565, n566, n567, n568, n569,
         n570, n571, n572, n573, n574, n575, n576, n577, n578, n579, n580,
         n581, n582, n583, n584, n585, n586, n587, n588, n589, n590, n591,
         n592, n593, n594, n595, n596, n597, n598, n599, n600, n601, n602,
         n603, n604, n605, n606, n607, n608, n609, n610, n611, n612, n613,
         n614, n615, n616, n617, n618, n619, n620, n621, n622, n623, n624,
         n625, n626, n627, n628, n629, n630, n631, n632, n633, n634, n635;
  wire   [10:0] addrD;
  wire   [15:0] addrT;
  wire   [1:0] \driver/start_history ;
  wire   [5:0] \decider/posy_m_obstacle_top ;
  wire   [15:0] \decider/obstacle_right ;
  wire   [7:3] \decider/posx_m_rex_left ;
  assign rw_o = \driver/*Logic0* ;

  DFFHQ \driver/en_o_reg  ( .D(\driver/N96 ), .CK(clk), .Q(en_o) );
  DFFHQ \driver/rst_o_reg  ( .D(n611), .CK(clk), .Q(rst_o) );
  EDFFHQ \driver/start_history_reg[0]  ( .D(start_i), .E(rstn), .CK(clk), .Q(
        \driver/start_history [0]) );
  EDFFHQ \driver/start_history_reg[1]  ( .D(\driver/start_history [0]), .E(
        rstn), .CK(clk), .Q(\driver/start_history [1]) );
  DFFHQ \driver/y_reg[5]  ( .D(n373), .CK(clk), .Q(addrD[5]) );
  DFFHQ \driver/y_reg[0]  ( .D(n372), .CK(clk), .Q(addrD[0]) );
  DFFHQ \driver/y_reg[1]  ( .D(n371), .CK(clk), .Q(addrD[1]) );
  DFFHQ \driver/y_reg[2]  ( .D(n370), .CK(clk), .Q(addrD[2]) );
  DFFHQ \driver/y_reg[3]  ( .D(n369), .CK(clk), .Q(addrD[3]) );
  DFFHQ \driver/y_reg[4]  ( .D(n368), .CK(clk), .Q(addrD[4]) );
  DFFHQ \driver/x_reg[4]  ( .D(n367), .CK(clk), .Q(addrD[10]) );
  DFFHQ \driver/x_reg[0]  ( .D(n366), .CK(clk), .Q(addrD[6]) );
  DFFHQ \driver/x_reg[1]  ( .D(n365), .CK(clk), .Q(addrD[7]) );
  DFFHQ \driver/x_reg[2]  ( .D(n364), .CK(clk), .Q(addrD[8]) );
  DFFHQ \driver/x_reg[3]  ( .D(n363), .CK(clk), .Q(addrD[9]) );
  DFFHQ \driver/state_reg[0]  ( .D(n361), .CK(clk), .Q(state[0]) );
  DFFHQ \driver/state_reg[1]  ( .D(n360), .CK(clk), .Q(state[1]) );
  DFFHQ \driver/state_reg[2]  ( .D(n362), .CK(clk), .Q(state[2]) );
  DFFHQ \driver/dori_o_reg  ( .D(n359), .CK(clk), .Q(dori_o) );
  DFFRHQ \decider/addrT_reg[0]  ( .D(n617), .CK(clk), .RN(rstn), .Q(addrT[0])
         );
  DFFRHQ \decider/addrT_reg[1]  ( .D(n618), .CK(clk), .RN(rstn), .Q(addrT[1])
         );
  DFFRHQ \decider/addrT_reg[2]  ( .D(n619), .CK(clk), .RN(rstn), .Q(addrT[2])
         );
  DFFRHQ \decider/addrT_reg[3]  ( .D(n620), .CK(clk), .RN(rstn), .Q(addrT[3])
         );
  DFFRHQ \decider/addrT_reg[4]  ( .D(n621), .CK(clk), .RN(rstn), .Q(addrT[4])
         );
  DFFRHQ \decider/addrT_reg[5]  ( .D(n622), .CK(clk), .RN(rstn), .Q(addrT[5])
         );
  DFFRHQ \decider/addrT_reg[6]  ( .D(n615), .CK(clk), .RN(rstn), .Q(addrT[6])
         );
  DFFRHQ \decider/addrT_reg[7]  ( .D(n614), .CK(clk), .RN(rstn), .Q(addrT[7])
         );
  DFFRHQ \decider/addrT_reg[8]  ( .D(n613), .CK(clk), .RN(rstn), .Q(addrT[8])
         );
  DFFRHQ \decider/addrT_reg[9]  ( .D(n612), .CK(clk), .RN(rstn), .Q(addrT[9])
         );
  DFFHQ \driver/db_o_reg[7]  ( .D(n610), .CK(clk), .Q(db_o[7]) );
  DFFHQ \driver/db_o_reg[0]  ( .D(n358), .CK(clk), .Q(db_o[0]) );
  DFFHQ \driver/db_o_reg[1]  ( .D(n357), .CK(clk), .Q(db_o[1]) );
  DFFHQ \driver/db_o_reg[2]  ( .D(n356), .CK(clk), .Q(db_o[2]) );
  DFFHQ \driver/db_o_reg[3]  ( .D(n355), .CK(clk), .Q(db_o[3]) );
  DFFHQ \driver/db_o_reg[4]  ( .D(n354), .CK(clk), .Q(db_o[4]) );
  DFFHQ \driver/db_o_reg[5]  ( .D(n353), .CK(clk), .Q(db_o[5]) );
  DFFHQ \driver/db_o_reg[6]  ( .D(n352), .CK(clk), .Q(db_o[6]) );
  ADDF \r50/U2_1  ( .A(\U3/U3/Z_1 ), .B(n627), .CI(\r50/carry[1] ), .CO(
        \r50/carry[2] ), .S(\decider/N88 ) );
  ADDF \r50/U2_2  ( .A(\U3/U3/Z_2 ), .B(n626), .CI(\r50/carry[2] ), .CO(
        \r50/carry[3] ), .S(\decider/N89 ) );
  ADDF \r50/U2_3  ( .A(\U3/U3/Z_3 ), .B(n625), .CI(\r50/carry[3] ), .CO(
        \r50/carry[4] ), .S(\decider/N90 ) );
  ADDF \r50/U2_4  ( .A(\U3/U3/Z_4 ), .B(n624), .CI(\r50/carry[4] ), .CO(
        \r50/carry[5] ), .S(\decider/N91 ) );
  ADDF \r50/U2_5  ( .A(\U3/U3/Z_5 ), .B(n623), .CI(\r50/carry[5] ), .CO(
        \r50/carry[6] ), .S(\decider/N92 ) );
  ADDF \r50/U2_6  ( .A(\U3/U3/Z_6 ), .B(n616), .CI(\r50/carry[6] ), .CO(
        \r50/carry[7] ), .S(\decider/N93 ) );
  ADDF \r50/U2_7  ( .A(\U3/U3/Z_7 ), .B(n616), .CI(\r50/carry[7] ), .CO(
        \r50/carry[8] ), .S(\decider/N94 ) );
  ADDF \r50/U2_8  ( .A(\U3/U3/Z_8 ), .B(n616), .CI(\r50/carry[8] ), .CO(
        \r50/carry[9] ), .S(\decider/N95 ) );
  ADDF \r50/U2_9  ( .A(\U3/U3/Z_9 ), .B(n616), .CI(\r50/carry[9] ), .S(
        \decider/N96 ) );
  ADDF \r61/S2_2_1  ( .A(\U3/U1/Z_2 ), .B(n393), .CI(\U3/U1/Z_1 ), .CO(
        \r61/CARRYB[2][1] ), .S(\r61/SUMB[2][1] ) );
  ADDF \r61/S1_2_0  ( .A(\r61/ab[2][0] ), .B(n392), .CI(\r61/SUMB[1][1] ), 
        .CO(\r61/CARRYB[2][0] ), .S(\decider/N57 ) );
  ADDF \r61/S2_3_2  ( .A(\U3/U1/Z_3 ), .B(n391), .CI(\U3/U1/Z_1 ), .CO(
        \r61/CARRYB[3][2] ), .S(\r61/SUMB[3][2] ) );
  ADDF \r61/S2_3_1  ( .A(\U3/U1/Z_3 ), .B(\r61/CARRYB[2][1] ), .CI(
        \r61/SUMB[2][2] ), .CO(\r61/CARRYB[3][1] ), .S(\r61/SUMB[3][1] ) );
  ADDF \r61/S1_3_0  ( .A(\r61/ab[3][0] ), .B(\r61/CARRYB[2][0] ), .CI(
        \r61/SUMB[2][1] ), .CO(\r61/CARRYB[3][0] ), .S(\decider/N58 ) );
  ADDF \r61/S2_4_2  ( .A(\U3/U1/Z_4 ), .B(\r61/CARRYB[3][2] ), .CI(\U3/U1/Z_2 ), .CO(\r61/CARRYB[4][2] ), .S(\r61/SUMB[4][2] ) );
  ADDF \r61/S2_4_1  ( .A(\U3/U1/Z_4 ), .B(\r61/CARRYB[3][1] ), .CI(
        \r61/SUMB[3][2] ), .CO(\r61/CARRYB[4][1] ), .S(\r61/SUMB[4][1] ) );
  ADDF \r61/S1_4_0  ( .A(\r61/ab[4][0] ), .B(\r61/CARRYB[3][0] ), .CI(
        \r61/SUMB[3][1] ), .CO(\r61/CARRYB[4][0] ), .S(\r61/PROD1[4] ) );
  ADDF \r61/S2_5_2  ( .A(\U3/U1/Z_8 ), .B(\r61/CARRYB[4][2] ), .CI(\U3/U1/Z_3 ), .CO(\r61/CARRYB[5][2] ), .S(\r61/SUMB[5][2] ) );
  ADDF \r61/S2_5_1  ( .A(\U3/U1/Z_8 ), .B(\r61/CARRYB[4][1] ), .CI(
        \r61/SUMB[4][2] ), .CO(\r61/CARRYB[5][1] ), .S(\r61/SUMB[5][1] ) );
  ADDF \r61/S2_6_2  ( .A(\U3/U1/Z_8 ), .B(\r61/CARRYB[5][2] ), .CI(\U3/U1/Z_4 ), .CO(\r61/SUMB[7][2] ), .S(\r61/SUMB[6][2] ) );
  ADDF \r61/S2_6_1  ( .A(\U3/U1/Z_8 ), .B(\r61/CARRYB[5][1] ), .CI(
        \r61/SUMB[5][2] ), .CO(\r61/CARRYB[6][1] ), .S(\r61/SUMB[6][1] ) );
  ADDF \r61/S2_7_1  ( .A(\U3/U1/Z_8 ), .B(\r61/CARRYB[6][1] ), .CI(
        \r61/SUMB[6][2] ), .CO(\r61/CARRYB[7][1] ), .S(\r61/SUMB[7][1] ) );
  ADDF \r61/S2_8_1  ( .A(\U3/U1/Z_8 ), .B(\r61/CARRYB[7][1] ), .CI(
        \r61/SUMB[7][2] ), .S(\r61/SUMB[8][1] ) );
  AND2 U302 ( .A(addrD[7]), .B(addrD[6]), .Y(n377) );
  AND2 U303 ( .A(addrD[8]), .B(n377), .Y(n378) );
  AND2 U304 ( .A(n383), .B(\r61/PROD1[4] ), .Y(n379) );
  AND2 U305 ( .A(n631), .B(n630), .Y(n380) );
  AND2 U306 ( .A(n632), .B(n631), .Y(n381) );
  AND2 U307 ( .A(n634), .B(\decider/sub_75/carry[4] ), .Y(n382) );
  AND2 U308 ( .A(\add_2_root_decider/add_109_3_cf/carry[3] ), .B(\decider/N58 ), .Y(n383) );
  AND2 U309 ( .A(\add_2_root_decider/add_109_3_cf/carry[7] ), .B(\decider/N62 ), .Y(n384) );
  AND2 U310 ( .A(\r61/CARRYB[4][0] ), .B(\r61/SUMB[4][1] ), .Y(n385) );
  AND2 U311 ( .A(n385), .B(\r61/SUMB[5][1] ), .Y(n386) );
  AND2 U312 ( .A(n386), .B(\r61/SUMB[6][1] ), .Y(n387) );
  AND2 U313 ( .A(addrD[9]), .B(n378), .Y(n388) );
  AND2 U314 ( .A(n384), .B(\decider/N63 ), .Y(n389) );
  AND2 U315 ( .A(n387), .B(\r61/SUMB[7][1] ), .Y(n390) );
  AND2 U316 ( .A(n405), .B(\U3/U1/Z_2 ), .Y(n391) );
  AND2 U317 ( .A(\r61/ab[1][0] ), .B(n405), .Y(n392) );
  AND2 U318 ( .A(n405), .B(\U3/U1/Z_1 ), .Y(n393) );
  INV U319 ( .A(n417), .Y(n394) );
  BUF U320 ( .I(n445), .O(n395) );
  BUF U321 ( .I(n446), .O(n396) );
  LOGIC_0 U322 ( .LOGIC_0_PIN(\driver/*Logic0* ) );
  NAND2 U323 ( .A(n397), .B(n398), .Y(\r50/carry[1] ) );
  XNOR2 U324 ( .A(n628), .B(\U3/U3/Z_0 ), .Y(\decider/N38 ) );
  INV U325 ( .A(n628), .Y(n397) );
  INV U326 ( .A(\U3/U3/Z_0 ), .Y(n398) );
  NAND2 U327 ( .A(n399), .B(n409), .Y(
        \add_2_root_decider/add_109_3_cf/carry[3] ) );
  XNOR2 U328 ( .A(\decider/N57 ), .B(
        \add_2_root_decider/add_109_3_cf/carry[2] ), .Y(\decider/N84 ) );
  INV U329 ( .A(\decider/N57 ), .Y(n399) );
  NAND2 U330 ( .A(n400), .B(n410), .Y(
        \add_2_root_decider/add_109_3_cf/carry[7] ) );
  XNOR2 U331 ( .A(\decider/N61 ), .B(
        \add_2_root_decider/add_109_3_cf/carry[6] ), .Y(\decider/N80 ) );
  INV U332 ( .A(\decider/N61 ), .Y(n400) );
  NAND2 U333 ( .A(addrD[3]), .B(n411), .Y(\sub_1_root_decider/sub_49/carry[4] ) );
  XNOR2 U334 ( .A(n633), .B(\sub_1_root_decider/sub_49/carry[3] ), .Y(
        \decider/posy_m_rex_top[3] ) );
  NAND2 U335 ( .A(addrD[5]), .B(n412), .Y(\sub_1_root_decider/sub_49/carry[6] ) );
  XNOR2 U336 ( .A(n629), .B(\sub_1_root_decider/sub_49/carry[5] ), .Y(
        \decider/posy_m_rex_top[5] ) );
  NAND2 U337 ( .A(n472), .B(n401), .Y(\decider/sub_45/carry[5] ) );
  XNOR2 U338 ( .A(addrD[10]), .B(\decider/sub_45/carry[4] ), .Y(
        \decider/posx_m_rex_left [7]) );
  INV U339 ( .A(\decider/sub_45/carry[4] ), .Y(n401) );
  NAND2 U340 ( .A(n402), .B(n403), .Y(\decider/sub_45/carry[4] ) );
  XNOR2 U341 ( .A(addrD[9]), .B(\decider/sub_45/carry[3] ), .Y(
        \decider/posx_m_rex_left [6]) );
  INV U342 ( .A(addrD[9]), .Y(n402) );
  INV U343 ( .A(\decider/sub_45/carry[3] ), .Y(n403) );
  NAND2 U344 ( .A(n476), .B(n404), .Y(\decider/sub_45/carry[3] ) );
  XNOR2 U345 ( .A(addrD[8]), .B(\decider/sub_45/carry[2] ), .Y(
        \decider/posx_m_rex_left [5]) );
  INV U346 ( .A(\decider/sub_45/carry[2] ), .Y(n404) );
  NAND2 U347 ( .A(n475), .B(n405), .Y(\decider/sub_45/carry[2] ) );
  XNOR2 U348 ( .A(addrD[7]), .B(addrD[6]), .Y(\decider/posx_m_rex_left [4]) );
  INV U349 ( .A(addrD[6]), .Y(n405) );
  NAND2 U350 ( .A(addrD[3]), .B(n406), .Y(\decider/sub_75/carry[4] ) );
  XNOR2 U351 ( .A(n633), .B(n381), .Y(\decider/posy_m_obstacle_top [3]) );
  INV U352 ( .A(n381), .Y(n406) );
  NAND2 U353 ( .A(addrD[5]), .B(n407), .Y(\decider/sub_75/carry[6] ) );
  XNOR2 U354 ( .A(n629), .B(n382), .Y(\decider/posy_m_obstacle_top [5]) );
  INV U355 ( .A(n382), .Y(n407) );
  XNOR2 U356 ( .A(n635), .B(\sub_0_root_decider/sub_73/carry[15] ), .Y(
        \decider/posx_m_obstacle_right[15] ) );
  NAND2 U357 ( .A(n402), .B(n413), .Y(\r180/carry[7] ) );
  XNOR2 U358 ( .A(addrD[9]), .B(n378), .Y(\decider/obstacle_right [6]) );
  NAND2 U359 ( .A(n472), .B(n408), .Y(\r180/carry[8] ) );
  XNOR2 U360 ( .A(addrD[10]), .B(\r180/carry[7] ), .Y(
        \decider/obstacle_right [7]) );
  INV U361 ( .A(\r180/carry[7] ), .Y(n408) );
  XOR2 U362 ( .A(addrD[7]), .B(addrD[6]), .Y(\driver/N44 ) );
  XOR2 U363 ( .A(addrD[8]), .B(n377), .Y(\driver/N45 ) );
  XOR2 U364 ( .A(addrD[9]), .B(n378), .Y(\driver/N46 ) );
  XOR2 U365 ( .A(addrD[10]), .B(n388), .Y(\driver/N47 ) );
  XOR2 U366 ( .A(\decider/N56 ), .B(\decider/N55 ), .Y(\decider/N85 ) );
  NAND2 U367 ( .A(\decider/N55 ), .B(\decider/N56 ), .Y(n409) );
  INV U368 ( .A(n409), .Y(\add_2_root_decider/add_109_3_cf/carry[2] ) );
  XOR2 U369 ( .A(\decider/N58 ), .B(\add_2_root_decider/add_109_3_cf/carry[3] ), .Y(\decider/N83 ) );
  XOR2 U370 ( .A(\r61/PROD1[4] ), .B(n383), .Y(\decider/N82 ) );
  XOR2 U371 ( .A(\decider/N60 ), .B(n379), .Y(\decider/N81 ) );
  NAND2 U372 ( .A(n379), .B(\decider/N60 ), .Y(n410) );
  INV U373 ( .A(n410), .Y(\add_2_root_decider/add_109_3_cf/carry[6] ) );
  XOR2 U374 ( .A(\decider/N62 ), .B(\add_2_root_decider/add_109_3_cf/carry[7] ), .Y(\decider/N79 ) );
  XOR2 U375 ( .A(\decider/N63 ), .B(n384), .Y(\decider/N78 ) );
  XOR2 U376 ( .A(\decider/N64 ), .B(n389), .Y(\decider/N77 ) );
  XOR2 U377 ( .A(\r61/ab[1][0] ), .B(n405), .Y(\decider/N56 ) );
  XOR2 U378 ( .A(\U3/U1/Z_1 ), .B(n405), .Y(\r61/SUMB[1][1] ) );
  XOR2 U379 ( .A(n631), .B(n630), .Y(\decider/posy_m_rex_top[1] ) );
  XOR2 U380 ( .A(n632), .B(n380), .Y(\decider/posy_m_rex_top[2] ) );
  NAND2 U381 ( .A(n632), .B(n380), .Y(n411) );
  INV U382 ( .A(n411), .Y(\sub_1_root_decider/sub_49/carry[3] ) );
  XOR2 U383 ( .A(n634), .B(\sub_1_root_decider/sub_49/carry[4] ), .Y(
        \decider/posy_m_rex_top[4] ) );
  NAND2 U384 ( .A(n634), .B(\sub_1_root_decider/sub_49/carry[4] ), .Y(n412) );
  INV U385 ( .A(n412), .Y(\sub_1_root_decider/sub_49/carry[5] ) );
  XOR2 U386 ( .A(n632), .B(n631), .Y(\decider/posy_m_obstacle_top [2]) );
  XOR2 U387 ( .A(n634), .B(\decider/sub_75/carry[4] ), .Y(
        \decider/posy_m_obstacle_top [4]) );
  XOR2 U388 ( .A(addrD[7]), .B(addrD[6]), .Y(\decider/obstacle_right [4]) );
  XOR2 U389 ( .A(addrD[8]), .B(n377), .Y(\decider/obstacle_right [5]) );
  NAND2 U390 ( .A(addrD[8]), .B(n377), .Y(n413) );
  XOR2 U391 ( .A(\U3/U1/Z_2 ), .B(n405), .Y(\r61/SUMB[2][2] ) );
  XOR2 U392 ( .A(\r61/CARRYB[4][0] ), .B(\r61/SUMB[4][1] ), .Y(\decider/N60 )
         );
  XOR2 U393 ( .A(n385), .B(\r61/SUMB[5][1] ), .Y(\decider/N61 ) );
  XOR2 U394 ( .A(n386), .B(\r61/SUMB[6][1] ), .Y(\decider/N62 ) );
  XOR2 U395 ( .A(n387), .B(\r61/SUMB[7][1] ), .Y(\decider/N63 ) );
  XOR2 U396 ( .A(n390), .B(\r61/SUMB[8][1] ), .Y(\decider/N64 ) );
  INV U397 ( .A(n414), .Y(\sub_0_root_decider/sub_73/carry[15] ) );
  NOR4BB U398 ( .AN(n415), .BN(\r180/carry[8] ), .C(
        \decider/obstacle_right [5]), .D(\decider/obstacle_right [4]), .Y(n414) );
  NOR2 U399 ( .A(\decider/obstacle_right [7]), .B(\decider/obstacle_right [6]), 
        .Y(n415) );
  OAI221 U400 ( .A0(n416), .A1(n417), .B0(n418), .B1(n419), .C0(n420), .Y(n610) );
  INV U401 ( .A(db_o[7]), .Y(n419) );
  AOI211 U402 ( .A0(n421), .A1(n422), .B0(n423), .C0(n424), .Y(n416) );
  INV U403 ( .A(n425), .Y(n424) );
  AOI32 U404 ( .A0(n426), .A1(n427), .A2(n428), .B0(n429), .B1(n430), .Y(n425)
         );
  OAI32 U405 ( .A0(addrT[1]), .A1(addrT[2]), .A2(n431), .B0(n427), .B1(n432), 
        .Y(n429) );
  OAI221 U406 ( .A0(addrT[4]), .A1(n433), .B0(n434), .B1(n435), .C0(n436), .Y(
        n423) );
  MX2 U407 ( .A(n437), .B(n438), .S0(addrT[3]), .Y(n436) );
  AOI2BB2 U408 ( .B0(n421), .B1(n439), .A0N(n432), .A1N(n440), .Y(n438) );
  INV U409 ( .A(n441), .Y(n437) );
  AOI221 U410 ( .A0(n442), .A1(n440), .B0(n443), .B1(addrT[5]), .C0(n444), .Y(
        n433) );
  MX2 U411 ( .A(addrT[3]), .B(addrT[6]), .S0(n426), .Y(n443) );
  MX2 U412 ( .A(\decider/N96 ), .B(addrT[9]), .S0(n395), .Y(n612) );
  MX2 U413 ( .A(\decider/N95 ), .B(addrT[8]), .S0(n395), .Y(n613) );
  MX2 U414 ( .A(\decider/N94 ), .B(addrT[7]), .S0(n395), .Y(n614) );
  MX2 U415 ( .A(\decider/N93 ), .B(addrT[6]), .S0(n395), .Y(n615) );
  NOR2B U416 ( .AN(\decider/sub_75/carry[6] ), .B(n396), .Y(n616) );
  MX2 U417 ( .A(\decider/N38 ), .B(addrT[0]), .S0(n395), .Y(n617) );
  MX2 U418 ( .A(\decider/N88 ), .B(addrT[1]), .S0(n395), .Y(n618) );
  MX2 U419 ( .A(\decider/N89 ), .B(addrT[2]), .S0(n395), .Y(n619) );
  MX2 U420 ( .A(\decider/N90 ), .B(addrT[3]), .S0(n395), .Y(n620) );
  MX2 U421 ( .A(\decider/N91 ), .B(addrT[4]), .S0(n395), .Y(n621) );
  MX2 U422 ( .A(\decider/N92 ), .B(addrT[5]), .S0(n395), .Y(n622) );
  AOI31 U423 ( .A0(\decider/posx_m_obstacle_right[15] ), .A1(n447), .A2(
        \r180/carry[8] ), .B0(n396), .Y(n445) );
  INV U424 ( .A(\decider/sub_75/carry[6] ), .Y(n447) );
  INV U425 ( .A(n448), .Y(n623) );
  MX2 U426 ( .A(\decider/posy_m_obstacle_top [5]), .B(
        \decider/posy_m_rex_top[5] ), .S0(n396), .Y(n448) );
  INV U427 ( .A(n449), .Y(n624) );
  MX2 U428 ( .A(\decider/posy_m_obstacle_top [4]), .B(
        \decider/posy_m_rex_top[4] ), .S0(n396), .Y(n449) );
  INV U429 ( .A(n450), .Y(n625) );
  MX2 U430 ( .A(\decider/posy_m_obstacle_top [3]), .B(
        \decider/posy_m_rex_top[3] ), .S0(n396), .Y(n450) );
  INV U431 ( .A(n451), .Y(n626) );
  MX2 U432 ( .A(\decider/posy_m_obstacle_top [2]), .B(
        \decider/posy_m_rex_top[2] ), .S0(n396), .Y(n451) );
  INV U433 ( .A(n452), .Y(n627) );
  MX2 U434 ( .A(addrD[1]), .B(\decider/posy_m_rex_top[1] ), .S0(n396), .Y(n452) );
  XOR2 U435 ( .A(addrD[0]), .B(n396), .Y(n628) );
  INV U436 ( .A(addrD[1]), .Y(n631) );
  MX2 U437 ( .A(n453), .B(n454), .S0(addrD[5]), .Y(n373) );
  OAI21 U438 ( .A0(addrD[4]), .A1(n455), .B0(n456), .Y(n454) );
  NOR2B U439 ( .AN(n457), .B(n455), .Y(n453) );
  MX2 U440 ( .A(n458), .B(n459), .S0(addrD[0]), .Y(n372) );
  MX2 U441 ( .A(n460), .B(n461), .S0(addrD[1]), .Y(n371) );
  INV U442 ( .A(n462), .Y(n461) );
  NOR2B U443 ( .AN(addrD[0]), .B(n455), .Y(n460) );
  MX2 U444 ( .A(n463), .B(n464), .S0(addrD[2]), .Y(n370) );
  OAI21 U445 ( .A0(addrD[1]), .A1(n455), .B0(n462), .Y(n464) );
  AOI2BB1 U446 ( .A0N(addrD[0]), .A1N(n455), .B0(n459), .Y(n462) );
  NOR3B U447 ( .AN(addrD[1]), .B(n455), .C(n630), .Y(n463) );
  MX2 U448 ( .A(n465), .B(n466), .S0(addrD[3]), .Y(n369) );
  NOR2B U449 ( .AN(n467), .B(n455), .Y(n465) );
  MX2 U450 ( .A(n468), .B(n469), .S0(addrD[4]), .Y(n368) );
  INV U451 ( .A(n456), .Y(n469) );
  AOI2BB1 U452 ( .A0N(addrD[3]), .A1N(n455), .B0(n466), .Y(n456) );
  OAI21 U453 ( .A0(n467), .A1(n455), .B0(n470), .Y(n466) );
  NOR3B U454 ( .AN(n467), .B(n455), .C(n633), .Y(n468) );
  OAI2BB2 U455 ( .B0(n471), .B1(n472), .A0N(\driver/N47 ), .A1N(n473), .Y(n367) );
  MX2 U456 ( .A(n473), .B(n474), .S0(addrD[6]), .Y(n366) );
  OAI2BB2 U457 ( .B0(n471), .B1(n475), .A0N(\driver/N44 ), .A1N(n473), .Y(n365) );
  OAI2BB2 U458 ( .B0(n471), .B1(n476), .A0N(\driver/N45 ), .A1N(n473), .Y(n364) );
  OAI2BB2 U459 ( .B0(n471), .B1(n402), .A0N(\driver/N46 ), .A1N(n473), .Y(n363) );
  NOR2B U460 ( .AN(n477), .B(n474), .Y(n473) );
  OAI21 U461 ( .A0(n478), .A1(n479), .B0(n480), .Y(n362) );
  NAND2 U462 ( .A(n481), .B(n480), .Y(n361) );
  MX2 U463 ( .A(n482), .B(n483), .S0(n484), .Y(n481) );
  AOI31 U464 ( .A0(cs_o[3]), .A1(addrD[8]), .A2(n485), .B0(n486), .Y(n482) );
  NOR3B U465 ( .AN(addrD[7]), .B(n405), .C(n487), .Y(n485) );
  NAND3 U466 ( .A(n488), .B(n480), .C(n489), .Y(n360) );
  MX2 U467 ( .A(n487), .B(n490), .S0(n484), .Y(n489) );
  OAI31 U468 ( .A0(n491), .A1(n611), .A2(n492), .B0(n479), .Y(n480) );
  INV U469 ( .A(n484), .Y(n479) );
  AOI211 U470 ( .A0(en_o), .A1(n491), .B0(n493), .C0(n471), .Y(n484) );
  INV U471 ( .A(n474), .Y(n471) );
  AOI31 U472 ( .A0(n494), .A1(addrD[5]), .A2(n457), .B0(n495), .Y(n474) );
  NOR3B U473 ( .AN(n467), .B(n633), .C(n634), .Y(n457) );
  NOR3B U474 ( .AN(addrD[1]), .B(n630), .C(n632), .Y(n467) );
  INV U475 ( .A(addrD[2]), .Y(n632) );
  INV U476 ( .A(addrD[0]), .Y(n630) );
  INV U477 ( .A(n496), .Y(n493) );
  NOR2B U478 ( .AN(n497), .B(n478), .Y(n491) );
  OAI2BB1 U479 ( .A0N(n498), .A1N(dori_o), .B0(n455), .Y(n359) );
  INV U480 ( .A(n458), .Y(n455) );
  NOR2B U481 ( .AN(n477), .B(n459), .Y(n458) );
  NOR2B U482 ( .AN(rstn), .B(n487), .Y(n477) );
  NOR2B U483 ( .AN(n496), .B(n470), .Y(n498) );
  INV U484 ( .A(n459), .Y(n470) );
  NOR2B U485 ( .AN(n499), .B(n495), .Y(n459) );
  OAI31 U486 ( .A0(n500), .A1(n488), .A2(n501), .B0(rstn), .Y(n495) );
  NAND2B U487 ( .AN(start_i), .B(en_o), .Y(n500) );
  OAI221 U488 ( .A0(n502), .A1(n503), .B0(n418), .B1(n504), .C0(n505), .Y(n358) );
  AOI222 U489 ( .A0(n506), .A1(addrD[0]), .B0(n507), .B1(n508), .C0(n509), 
        .C1(addrD[6]), .Y(n505) );
  OAI211 U490 ( .A0(n510), .A1(n511), .B0(n512), .C0(n513), .Y(n508) );
  AOI221 U491 ( .A0(n514), .A1(n515), .B0(n516), .B1(n517), .C0(n442), .Y(n513) );
  NOR2B U492 ( .AN(n518), .B(addrT[3]), .Y(n516) );
  INV U493 ( .A(n519), .Y(n511) );
  AOI2BB1 U494 ( .A0N(n427), .A1N(n520), .B0(n521), .Y(n510) );
  INV U495 ( .A(db_o[0]), .Y(n504) );
  OAI211 U496 ( .A0(n475), .A1(n420), .B0(n522), .C0(n523), .Y(n357) );
  AOI222 U497 ( .A0(db_o[1]), .A1(n524), .B0(n507), .B1(n525), .C0(n506), .C1(
        addrD[1]), .Y(n523) );
  OAI211 U498 ( .A0(n526), .A1(n440), .B0(n527), .C0(n528), .Y(n525) );
  NOR2B U499 ( .AN(n512), .B(n529), .Y(n528) );
  MX2 U500 ( .A(n530), .B(n442), .S0(addrT[1]), .Y(n529) );
  NOR2B U501 ( .AN(n434), .B(n435), .Y(n530) );
  INV U502 ( .A(n531), .Y(n512) );
  OAI33 U503 ( .A0(n532), .A1(n533), .A2(n431), .B0(n534), .B1(addrT[4]), .B2(
        n535), .Y(n531) );
  NOR2 U504 ( .A(n520), .B(n422), .Y(n535) );
  NOR2B U505 ( .AN(n521), .B(n536), .Y(n422) );
  AOI2BB1 U506 ( .A0N(n515), .A1N(n537), .B0(n538), .Y(n533) );
  AOI33 U507 ( .A0(n430), .A1(n439), .A2(n517), .B0(n539), .B1(addrT[0]), .B2(
        n519), .Y(n527) );
  NOR3B U508 ( .AN(n537), .B(addrT[1]), .C(addrT[6]), .Y(n519) );
  AOI31 U509 ( .A0(n540), .A1(n537), .A2(addrT[3]), .B0(n541), .Y(n526) );
  AOI31 U510 ( .A0(n539), .A1(n515), .A2(n542), .B0(n543), .Y(n522) );
  INV U511 ( .A(addrD[7]), .Y(n475) );
  NAND2B U512 ( .AN(n544), .B(n545), .Y(n356) );
  AOI222 U513 ( .A0(db_o[2]), .A1(n524), .B0(n507), .B1(n546), .C0(n506), .C1(
        addrD[2]), .Y(n545) );
  INV U514 ( .A(n547), .Y(n546) );
  AOI221 U515 ( .A0(n548), .A1(addrT[0]), .B0(n536), .B1(n549), .C0(n550), .Y(
        n547) );
  INV U516 ( .A(n551), .Y(n548) );
  AOI31 U517 ( .A0(addrT[2]), .A1(n515), .A2(n552), .B0(n442), .Y(n551) );
  OAI221 U518 ( .A0(n553), .A1(n554), .B0(n476), .B1(n420), .C0(n555), .Y(n544) );
  INV U519 ( .A(addrD[8]), .Y(n476) );
  NOR2B U520 ( .AN(n520), .B(n440), .Y(n553) );
  NOR2B U521 ( .AN(n434), .B(n532), .Y(n520) );
  INV U522 ( .A(n556), .Y(n355) );
  AOI211 U523 ( .A0(db_o[3]), .A1(n524), .B0(n557), .C0(n558), .Y(n556) );
  OAI222 U524 ( .A0(n559), .A1(n417), .B0(n560), .B1(n554), .C0(n633), .C1(
        n561), .Y(n557) );
  INV U525 ( .A(addrD[3]), .Y(n633) );
  NOR2B U526 ( .AN(n539), .B(addrT[0]), .Y(n560) );
  AOI211 U527 ( .A0(n549), .A1(n562), .B0(n550), .C0(n444), .Y(n559) );
  OAI211 U528 ( .A0(n515), .A1(n563), .B0(n435), .C0(n564), .Y(n550) );
  INV U529 ( .A(n541), .Y(n435) );
  INV U530 ( .A(n565), .Y(n354) );
  AOI211 U531 ( .A0(db_o[4]), .A1(n524), .B0(n566), .C0(n558), .Y(n565) );
  OAI222 U532 ( .A0(n567), .A1(n554), .B0(n568), .B1(n417), .C0(n634), .C1(
        n561), .Y(n566) );
  INV U533 ( .A(addrD[4]), .Y(n634) );
  AOI211 U534 ( .A0(n441), .A1(n532), .B0(n569), .C0(n570), .Y(n568) );
  OAI31 U535 ( .A0(n571), .A1(n515), .A2(n534), .B0(n572), .Y(n569) );
  NOR2 U536 ( .A(n541), .B(n549), .Y(n572) );
  NOR2B U537 ( .AN(n552), .B(addrT[2]), .Y(n549) );
  NOR2B U538 ( .AN(n552), .B(addrT[3]), .Y(n541) );
  MX2 U539 ( .A(n573), .B(n574), .S0(addrT[1]), .Y(n441) );
  NOR2B U540 ( .AN(n575), .B(n434), .Y(n573) );
  AOI2BB1 U541 ( .A0N(n427), .A1N(n571), .B0(n576), .Y(n567) );
  MX2 U542 ( .A(n518), .B(addrT[1]), .S0(addrT[3]), .Y(n576) );
  INV U543 ( .A(n426), .Y(n518) );
  INV U544 ( .A(n577), .Y(n353) );
  AOI211 U545 ( .A0(db_o[5]), .A1(n524), .B0(n578), .C0(n558), .Y(n577) );
  NAND2 U546 ( .A(n420), .B(n555), .Y(n558) );
  INV U547 ( .A(n543), .Y(n555) );
  NOR2B U548 ( .AN(n579), .B(n502), .Y(n543) );
  OAI31 U549 ( .A0(n501), .A1(start_i), .A2(n488), .B0(n503), .Y(n579) );
  INV U550 ( .A(n492), .Y(n503) );
  INV U551 ( .A(n580), .Y(n488) );
  INV U552 ( .A(\driver/start_history [1]), .Y(n501) );
  INV U553 ( .A(n509), .Y(n420) );
  NOR2B U554 ( .AN(n581), .B(n502), .Y(n509) );
  OAI222 U555 ( .A0(n582), .A1(n554), .B0(n583), .B1(n417), .C0(n629), .C1(
        n561), .Y(n578) );
  INV U556 ( .A(addrD[5]), .Y(n629) );
  NOR2B U557 ( .AN(n584), .B(n570), .Y(n583) );
  OAI211 U558 ( .A0(n563), .A1(n562), .B0(n564), .C0(n585), .Y(n570) );
  AOI31 U559 ( .A0(n427), .A1(n532), .A2(n575), .B0(n444), .Y(n585) );
  AOI31 U560 ( .A0(n586), .A1(n439), .A2(addrT[5]), .B0(n421), .Y(n564) );
  NOR2B U561 ( .AN(n587), .B(n588), .Y(n421) );
  NOR2B U562 ( .AN(n537), .B(addrT[3]), .Y(n586) );
  INV U563 ( .A(n514), .Y(n563) );
  NOR2B U564 ( .AN(n539), .B(addrT[5]), .Y(n514) );
  AOI211 U565 ( .A0(n538), .A1(addrT[3]), .B0(n539), .C0(n536), .Y(n582) );
  INV U566 ( .A(n589), .Y(n352) );
  AOI221 U567 ( .A0(n394), .A1(n590), .B0(db_o[6]), .B1(n524), .C0(n591), .Y(
        n589) );
  OAI31 U568 ( .A0(n554), .A1(n538), .A2(n571), .B0(n561), .Y(n591) );
  INV U569 ( .A(n506), .Y(n561) );
  NOR2B U570 ( .AN(n486), .B(n502), .Y(n506) );
  INV U571 ( .A(n592), .Y(n502) );
  INV U572 ( .A(n539), .Y(n571) );
  INV U573 ( .A(n542), .Y(n554) );
  NOR2B U574 ( .AN(n587), .B(n417), .Y(n542) );
  INV U575 ( .A(n507), .Y(n417) );
  NOR2 U576 ( .A(n537), .B(addrT[5]), .Y(n587) );
  INV U577 ( .A(n418), .Y(n524) );
  OAI221 U578 ( .A0(n593), .A1(n515), .B0(n432), .B1(n440), .C0(n594), .Y(n590) );
  NOR2B U579 ( .AN(n584), .B(n595), .Y(n594) );
  MX2 U580 ( .A(n596), .B(n597), .S0(addrT[4]), .Y(n595) );
  AOI211 U581 ( .A0(n562), .A1(n440), .B0(n532), .C0(n431), .Y(n597) );
  INV U582 ( .A(n538), .Y(n562) );
  NOR2B U583 ( .AN(addrT[0]), .B(n515), .Y(n538) );
  OAI2BB1 U584 ( .A0N(addrT[5]), .A1N(n598), .B0(n599), .Y(n596) );
  INV U585 ( .A(n444), .Y(n599) );
  NOR3B U586 ( .AN(n521), .B(n440), .C(n534), .Y(n444) );
  INV U587 ( .A(n540), .Y(n534) );
  NOR2B U588 ( .AN(addrT[6]), .B(addrT[5]), .Y(n540) );
  NOR2B U589 ( .AN(addrT[2]), .B(addrT[3]), .Y(n521) );
  MX2 U590 ( .A(n439), .B(n426), .S0(n532), .Y(n598) );
  NAND2B U591 ( .AN(n427), .B(n426), .Y(n439) );
  NOR2B U592 ( .AN(addrT[2]), .B(n515), .Y(n426) );
  AOI221 U593 ( .A0(n575), .A1(n600), .B0(n434), .B1(n428), .C0(n552), .Y(n584) );
  NOR2B U594 ( .AN(n575), .B(addrT[4]), .Y(n552) );
  NOR2B U595 ( .AN(n532), .B(addrT[1]), .Y(n600) );
  INV U596 ( .A(n536), .Y(n440) );
  NOR2B U597 ( .AN(n515), .B(addrT[0]), .Y(n536) );
  INV U598 ( .A(n574), .Y(n432) );
  NOR2B U599 ( .AN(n575), .B(addrT[2]), .Y(n574) );
  NOR2B U600 ( .AN(addrT[5]), .B(addrT[6]), .Y(n575) );
  INV U601 ( .A(addrT[1]), .Y(n515) );
  AOI21 U602 ( .A0(n427), .A1(n428), .B0(n442), .Y(n593) );
  NOR2B U603 ( .AN(n539), .B(n431), .Y(n442) );
  INV U604 ( .A(n517), .Y(n431) );
  NOR2B U605 ( .AN(n588), .B(addrT[5]), .Y(n517) );
  INV U606 ( .A(addrT[6]), .Y(n588) );
  NOR2B U607 ( .AN(addrT[3]), .B(n434), .Y(n539) );
  INV U608 ( .A(addrT[2]), .Y(n434) );
  NOR2B U609 ( .AN(n430), .B(addrT[6]), .Y(n428) );
  NOR2B U610 ( .AN(n532), .B(n537), .Y(n430) );
  INV U611 ( .A(addrT[4]), .Y(n537) );
  INV U612 ( .A(addrT[3]), .Y(n532) );
  INV U613 ( .A(addrT[0]), .Y(n427) );
  NOR4 U614 ( .A(addrT[9]), .B(addrT[8]), .C(addrT[7]), .D(n601), .Y(n507) );
  OAI211 U615 ( .A0(n602), .A1(n396), .B0(n603), .C0(n592), .Y(n601) );
  NOR2B U616 ( .AN(n418), .B(n611), .Y(n592) );
  INV U617 ( .A(rstn), .Y(n611) );
  OAI211 U618 ( .A0(n604), .A1(\driver/N96 ), .B0(n496), .C0(n499), .Y(n418)
         );
  INV U619 ( .A(n494), .Y(n499) );
  NOR2B U620 ( .AN(en_o), .B(n487), .Y(n494) );
  INV U621 ( .A(n603), .Y(n487) );
  OAI31 U622 ( .A0(n492), .A1(n581), .A2(n486), .B0(en_o), .Y(n496) );
  NOR3B U623 ( .AN(n483), .B(state[2]), .C(n490), .Y(n486) );
  NOR3B U624 ( .AN(n490), .B(state[2]), .C(n483), .Y(n581) );
  INV U625 ( .A(state[1]), .Y(n490) );
  NOR2B U626 ( .AN(n478), .B(n497), .Y(n492) );
  INV U627 ( .A(state[2]), .Y(n478) );
  NOR2B U628 ( .AN(rstn), .B(n580), .Y(n604) );
  NOR2B U629 ( .AN(state[2]), .B(n497), .Y(n580) );
  NAND2 U630 ( .A(state[0]), .B(state[1]), .Y(n497) );
  NOR3B U631 ( .AN(n483), .B(state[2]), .C(state[1]), .Y(n603) );
  INV U632 ( .A(state[0]), .Y(n483) );
  NOR3B U633 ( .AN(\decider/posx_m_obstacle_right[15] ), .B(n635), .C(
        \decider/sub_75/carry[6] ), .Y(n602) );
  NOR2B U634 ( .AN(rstn), .B(en_o), .Y(\driver/N96 ) );
  NOR2B U635 ( .AN(n396), .B(addrD[6]), .Y(\decider/N55 ) );
  NOR2B U636 ( .AN(addrD[10]), .B(n402), .Y(cs_o[3]) );
  NOR2B U637 ( .AN(addrD[10]), .B(addrD[9]), .Y(cs_o[2]) );
  NOR2B U638 ( .AN(n472), .B(n402), .Y(cs_o[1]) );
  MX2 U639 ( .A(\decider/N77 ), .B(\decider/N64 ), .S0(n396), .Y(\U3/U3/Z_9 )
         );
  MX2 U640 ( .A(\decider/N78 ), .B(\decider/N63 ), .S0(n396), .Y(\U3/U3/Z_8 )
         );
  MX2 U641 ( .A(\decider/N79 ), .B(\decider/N62 ), .S0(n396), .Y(\U3/U3/Z_7 )
         );
  MX2 U642 ( .A(\decider/N80 ), .B(\decider/N61 ), .S0(n396), .Y(\U3/U3/Z_6 )
         );
  MX2 U643 ( .A(\decider/N81 ), .B(\decider/N60 ), .S0(n396), .Y(\U3/U3/Z_5 )
         );
  MX2 U644 ( .A(\decider/N82 ), .B(\r61/PROD1[4] ), .S0(n396), .Y(\U3/U3/Z_4 )
         );
  MX2 U645 ( .A(\decider/N83 ), .B(\decider/N58 ), .S0(n396), .Y(\U3/U3/Z_3 )
         );
  MX2 U646 ( .A(\decider/N84 ), .B(\decider/N57 ), .S0(n396), .Y(\U3/U3/Z_2 )
         );
  MX2 U647 ( .A(\decider/N85 ), .B(\decider/N56 ), .S0(n446), .Y(\U3/U3/Z_1 )
         );
  NAND2 U648 ( .A(addrD[6]), .B(n396), .Y(\U3/U3/Z_0 ) );
  NOR2B U649 ( .AN(n635), .B(n396), .Y(\U3/U1/Z_8 ) );
  INV U650 ( .A(\r180/carry[8] ), .Y(n635) );
  OAI2BB1 U651 ( .A0N(n605), .A1N(\decider/obstacle_right [7]), .B0(n606), .Y(
        \U3/U1/Z_4 ) );
  INV U652 ( .A(\r61/ab[4][0] ), .Y(n606) );
  NOR2B U653 ( .AN(\decider/posx_m_rex_left [7]), .B(n605), .Y(\r61/ab[4][0] )
         );
  OAI2BB1 U654 ( .A0N(n605), .A1N(\decider/obstacle_right [6]), .B0(n607), .Y(
        \U3/U1/Z_3 ) );
  INV U655 ( .A(\r61/ab[3][0] ), .Y(n607) );
  NOR2B U656 ( .AN(\decider/posx_m_rex_left [6]), .B(n605), .Y(\r61/ab[3][0] )
         );
  OAI2BB1 U657 ( .A0N(n605), .A1N(\decider/obstacle_right [5]), .B0(n608), .Y(
        \U3/U1/Z_2 ) );
  INV U658 ( .A(\r61/ab[2][0] ), .Y(n608) );
  NOR2B U659 ( .AN(\decider/posx_m_rex_left [5]), .B(n605), .Y(\r61/ab[2][0] )
         );
  OAI2BB1 U660 ( .A0N(n605), .A1N(\decider/obstacle_right [4]), .B0(n609), .Y(
        \U3/U1/Z_1 ) );
  INV U661 ( .A(\r61/ab[1][0] ), .Y(n609) );
  NOR2B U662 ( .AN(\decider/posx_m_rex_left [4]), .B(n605), .Y(\r61/ab[1][0] )
         );
  INV U663 ( .A(n396), .Y(n605) );
  NOR4BB U664 ( .AN(\decider/sub_45/carry[5] ), .BN(cs_o[0]), .C(addrD[8]), 
        .D(\sub_1_root_decider/sub_49/carry[6] ), .Y(n446) );
  NOR2B U665 ( .AN(n472), .B(addrD[9]), .Y(cs_o[0]) );
  INV U666 ( .A(addrD[10]), .Y(n472) );
endmodule

