
module FDE_Rex_Runner ( clk, rstn, jmp_key, db_o, dori_o, cs_o, en_o, rw_o, 
        rst_o, state );
  output [7:0] db_o;
  output [3:0] cs_o;
  output [2:0] state;
  input clk, rstn, jmp_key;
  output dori_o, en_o, rw_o, rst_o;
  wire   start, \driver/N96 , \driver/N47 , \driver/N46 , \driver/N45 ,
         \driver/N44 , \driver/N17 , \decider/N102 , \decider/N101 ,
         \decider/N100 , \decider/N99 , \decider/N98 , \decider/N97 ,
         \decider/N96 , \decider/N95 , \decider/N94 , \decider/N93 ,
         \decider/N92 , \decider/N91 , \decider/N90 , \decider/N89 ,
         \decider/N88 , \decider/N87 , \decider/N86 , \decider/N85 ,
         \decider/N84 , \decider/N83 , \decider/N82 , \decider/N81 ,
         \decider/N80 , \decider/N79 , \decider/N78 , \decider/N77 ,
         \decider/N76 , \decider/N75 , \decider/N74 , \decider/N73 ,
         \decider/N72 , \decider/N71 , \decider/N65 , \decider/N64 ,
         \decider/N63 , \decider/N62 , \decider/N61 , \decider/N60 ,
         \decider/N58 , \decider/N57 , \decider/posy_m_rex_top[1] ,
         \decider/posy_m_rex_top[2] , \decider/posy_m_rex_top[3] ,
         \decider/posy_m_rex_top[4] , \decider/posy_m_rex_top[5] ,
         \decider/posy_m_rex_top[6] , \decider/posy_m_rex_top[7] ,
         \decider/posy_m_rex_top[8] , \decider/posy_m_rex_top[9] ,
         \decider/posy_m_rex_top[10] , \decider/posy_m_rex_top[11] ,
         \decider/posy_m_rex_top[12] , \decider/posy_m_rex_top[13] ,
         \decider/posy_m_rex_top[14] , \decider/posy_m_rex_top[15] ,
         \clock_divider/N30 , \clock_divider/N29 , \clock_divider/N28 ,
         \clock_divider/N27 , \clock_divider/N26 , \clock_divider/N25 ,
         \clock_divider/N24 , \clock_divider/N23 , \clock_divider/N22 ,
         \clock_divider/N21 , \clock_divider/N20 , \clock_divider/N19 ,
         \clock_divider/N18 , \clock_divider/N17 , \clock_divider/N16 ,
         \clock_divider/N15 , \clock_divider/N14 , \clock_divider/N13 ,
         \clock_divider/N12 , \clock_divider/N11 , \clock_divider/N10 ,
         \clock_divider/N9 , \clock_divider/N8 , \clock_divider/N7 ,
         \clock_divider/N6 , \clock_divider/cnt5k[0] ,
         \clock_divider/cnt5k[1] , \clock_divider/cnt5k[2] ,
         \clock_divider/cnt5k[3] , \clock_divider/cnt5k[4] ,
         \clock_divider/cnt5k[5] , \clock_divider/cnt5k[6] ,
         \clock_divider/cnt5k[7] , \clock_divider/cnt5k[8] ,
         \clock_divider/cnt5k[9] , \clock_divider/cnt5k[10] ,
         \clock_divider/cnt5k[11] , \clock_divider/cnt5k[12] , \U1/U2/Z_0 ,
         \U1/U2/Z_1 , \U1/U2/Z_2 , \U1/U2/Z_3 , \U1/U2/Z_4 , \U1/U2/Z_5 ,
         \U1/U2/Z_6 , \U1/U2/Z_7 , \U1/U2/Z_8 , \U1/U2/Z_9 , \U1/U2/Z_10 ,
         \U1/U2/Z_11 , \U1/U2/Z_12 , \U1/U2/Z_13 , \U1/U2/Z_14 , \U1/U2/Z_15 ,
         \U1/U3/Z_0 , \U1/U3/Z_1 , \U1/U3/Z_2 , \U1/U3/Z_3 , \U1/U3/Z_4 ,
         \U1/U5/Z_0 , \U1/U5/Z_1 , \U1/U5/Z_2 , \U1/U5/Z_3 , \U1/U5/Z_4 ,
         \U1/U5/Z_5 , \U1/U5/Z_6 , \U1/U5/Z_7 , \U1/U5/Z_8 , \U1/U5/Z_9 ,
         \U1/U5/Z_10 , \U1/U5/Z_11 , \U1/U5/Z_12 , \U1/U5/Z_13 , \U1/U5/Z_14 ,
         \U1/U5/Z_15 , n356, n366, n367, n368, n369, n370, n371, n372, n375,
         n376, n377, n378, n379, n380, n381, n382, n383, n384, n385, n386,
         n387, n388, n389, n390, n391, n392, n393, n394, n395, n396, n397,
         n398, \decider/sub_75/carry[6] , \decider/sub_75/carry[5] ,
         \sub_0_root_decider/sub_73/carry[15] ,
         \sub_0_root_decider/sub_49/carry[2] ,
         \sub_0_root_decider/sub_49/carry[3] ,
         \sub_0_root_decider/sub_49/carry[5] ,
         \sub_0_root_decider/sub_49/carry[6] ,
         \sub_0_root_decider/sub_49/carry[7] ,
         \sub_0_root_decider/sub_49/carry[8] ,
         \sub_0_root_decider/sub_49/carry[9] ,
         \sub_0_root_decider/sub_49/carry[10] ,
         \sub_0_root_decider/sub_49/carry[11] ,
         \sub_0_root_decider/sub_49/carry[12] ,
         \sub_0_root_decider/sub_49/carry[13] ,
         \sub_0_root_decider/sub_49/carry[14] ,
         \sub_0_root_decider/sub_49/carry[15] , \r250/carry[15] ,
         \r250/carry[14] , \r250/carry[13] , \r250/carry[12] ,
         \r250/carry[11] , \r250/carry[10] , \r250/carry[9] , \r250/carry[8] ,
         \r250/carry[7] , \r250/carry[6] , \r250/carry[5] , \r250/carry[4] ,
         \r250/carry[3] , \r250/carry[2] , \r250/carry[1] , \r191/B_not[15] ,
         \r191/B_not[14] , \r191/B_not[13] , \r191/B_not[12] ,
         \r191/B_not[11] , \r191/B_not[10] , \r191/B_not[9] , \r191/B_not[8] ,
         \r191/B_not[7] , \r191/B_not[6] , \r191/B_not[5] , \r191/B_not[4] ,
         \r191/B_not[3] , \r191/carry[15] , \r191/carry[14] , \r191/carry[13] ,
         \r191/carry[12] , \r191/carry[11] , \r191/carry[10] , \r191/carry[9] ,
         \r191/carry[8] , \r191/carry[7] , \r191/carry[6] , \r191/carry[5] ,
         \r191/carry[4] , \r191/carry[3] , \r187/B_not[15] , \r187/B_not[14] ,
         \r187/B_not[13] , \r187/B_not[12] , \r187/B_not[11] ,
         \r187/B_not[10] , \r187/B_not[9] , \r187/B_not[8] , \r187/B_not[7] ,
         \r187/B_not[6] , \r187/B_not[5] , \r187/B_not[4] , \r187/B_not[3] ,
         \r187/B_not[2] , \r187/B_not[1] , \r187/B_not[0] , \r187/carry[15] ,
         \r187/carry[14] , \r187/carry[13] , \r187/carry[12] ,
         \r187/carry[11] , \r187/carry[10] , \r187/carry[9] , \r187/carry[8] ,
         \r187/carry[7] , \r187/carry[6] , \r187/carry[5] , \r187/carry[4] ,
         \r187/carry[3] , \r187/carry[2] , \r187/carry[1] , \driver/*Logic0* ,
         \r62/A1[9] , \r62/A1[11] , \r62/A1[13] , \r62/PROD1[4] ,
         \r62/SUMB[1][2] , \r62/SUMB[1][3] , \r62/SUMB[2][2] ,
         \r62/SUMB[2][3] , \r62/SUMB[3][2] , \r62/SUMB[3][3] ,
         \r62/SUMB[4][2] , \r62/SUMB[4][3] , \r62/SUMB[5][2] ,
         \r62/SUMB[5][3] , \r62/SUMB[6][2] , \r62/SUMB[6][3] ,
         \r62/SUMB[7][2] , \r62/SUMB[7][3] , \r62/SUMB[8][2] ,
         \r62/SUMB[8][3] , \r62/SUMB[9][2] , \r62/SUMB[9][3] ,
         \r62/SUMB[10][2] , \r62/SUMB[10][3] , \r62/SUMB[11][2] ,
         \r62/SUMB[11][3] , \r62/SUMB[12][0] , \r62/SUMB[12][2] ,
         \r62/SUMB[12][3] , \r62/CARRYB[2][2] , \r62/CARRYB[2][3] ,
         \r62/CARRYB[3][0] , \r62/CARRYB[3][2] , \r62/CARRYB[3][3] ,
         \r62/CARRYB[4][0] , \r62/CARRYB[4][2] , \r62/CARRYB[4][3] ,
         \r62/CARRYB[5][2] , \r62/CARRYB[5][3] , \r62/CARRYB[6][2] ,
         \r62/CARRYB[6][3] , \r62/CARRYB[7][2] , \r62/CARRYB[7][3] ,
         \r62/CARRYB[8][2] , \r62/CARRYB[8][3] , \r62/CARRYB[9][2] ,
         \r62/CARRYB[9][3] , \r62/CARRYB[10][2] , \r62/CARRYB[10][3] ,
         \r62/CARRYB[11][2] , \r62/CARRYB[11][3] , \r62/CARRYB[12][2] ,
         \r62/ab[0][2] , \r62/ab[1][2] , \r62/ab[2][0] , \r62/ab[2][2] ,
         \r62/ab[3][0] , \r62/ab[3][2] , \r62/ab[4][0] , \r62/ab[4][2] ,
         \r62/ab[5][2] , \r62/ab[6][2] , \r62/ab[7][2] , \r62/ab[8][2] ,
         \r62/ab[9][2] , \r62/ab[10][2] , \r62/ab[11][2] , \r62/ab[12][2] ,
         \decider/sub_45/carry[2] , \decider/sub_45/carry[3] ,
         \decider/sub_45/carry[4] , \decider/sub_45/carry[5] , \r50/carry[7] ,
         \r50/carry[4] , \r50/carry[2] , n402, n403, n404, n405, n406, n407,
         n408, n409, n410, n411, n412, n413, n414, n415, n416, n417, n418,
         n419, n420, n421, n422, n423, n424, n425, n426, n427, n428, n429,
         n430, n431, n432, n433, n434, n435, n436, n437, n438, n439, n440,
         n441, n442, n443, n444, n445, n446, n447, n448, n449, n450, n451,
         n452, n453, n454, n455, n456, n457, n458, n459, n460, n461, n462,
         n463, n464, n465, n466, n467, n468, n469, n470, n471, n472, n473,
         n474, n475, n476, n477, n478, n479, n480, n481, n482, n483, n484,
         n485, n486, n487, n488, n489, n490, n491, n492, n493, n494, n495,
         n496, n497, n498, n499, n500, n501, n502, n503, n504, n505, n506,
         n507, n508, n509, n510, n511, n512, n513, n514, n515, n516, n517,
         n518, n519, n520, n521, n522, n523, n524, n525, n526, n527, n528,
         n529, n530, n531, n532, n533, n534, n535, n536, n537, n538, n539,
         n540, n541, n542, n543, n544, n545, n546, n547, n548, n549, n550,
         n551, n552, n553, n554, n555, n556, n557, n558, n559, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n570, n571, n572,
         n573, n574, n575, n576, n577, n578, n579, n580, n581, n582, n583,
         n584, n585, n586, n587, n588, n589, n590, n591, n592, n593, n594,
         n595, n596, n597, n598, n599, n600, n601, n602, n603, n604, n605,
         n606, n607, n608, n609, n610, n611, n612, n613, n614, n615, n616,
         n617, n618, n619, n620, n621, n622, n623, n624, n625, n626, n627,
         n628, n629, n630, n631, n632, n633, n634, n635, n636, n637, n638,
         n639, n640, n641, n642, n643, n644, n645, n646, n647, n648, n649,
         n650, n651, n652, n653, n654, n655, n656, n657, n658, n659, n660,
         n661, n662, n663, n664, n665, n666, n667, n668, n669, n670, n671,
         n672, n673, n674, n675, n676, n677, n678, n679, n680, n681, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736;
  wire   [10:0] addrD;
  wire   [15:0] addrT;
  wire   [1:0] \driver/start_history ;
  wire   [5:0] \decider/posy_m_obstacle_top ;
  wire   [15:0] \decider/obstacle_right ;
  wire   [7:3] \decider/posx_m_rex_left ;
  wire   [15:0] \decider/rex_top ;
  tri   clk;
  tri   rstn;
  tri   jmp_key;
  tri   [15:0] rex_down;
  tri   [15:0] obstacle_left;
  assign rw_o = \driver/*Logic0* ;

  DFFHQ \driver/en_o_reg  ( .D(\driver/N96 ), .CK(clk), .Q(en_o) );
  DFFHQ \driver/rst_o_reg  ( .D(\driver/N17 ), .CK(clk), .Q(rst_o) );
  DFFRHQ \clock_divider/cnt5k_reg[12]  ( .D(\clock_divider/N30 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[12] ) );
  DFFRHQ \clock_divider/clk_12Hz_reg  ( .D(n356), .CK(clk), .RN(rstn), .Q(
        start) );
  EDFFHQ \driver/start_history_reg[0]  ( .D(start), .E(rstn), .CK(clk), .Q(
        \driver/start_history [0]) );
  EDFFHQ \driver/start_history_reg[1]  ( .D(\driver/start_history [0]), .E(
        rstn), .CK(clk), .Q(\driver/start_history [1]) );
  DFFHQ \driver/y_reg[5]  ( .D(n398), .CK(clk), .Q(addrD[5]) );
  DFFHQ \driver/y_reg[0]  ( .D(n397), .CK(clk), .Q(addrD[0]) );
  DFFHQ \driver/y_reg[1]  ( .D(n396), .CK(clk), .Q(addrD[1]) );
  DFFHQ \driver/y_reg[2]  ( .D(n395), .CK(clk), .Q(addrD[2]) );
  DFFHQ \driver/y_reg[3]  ( .D(n394), .CK(clk), .Q(addrD[3]) );
  DFFHQ \driver/y_reg[4]  ( .D(n393), .CK(clk), .Q(addrD[4]) );
  DFFHQ \driver/x_reg[4]  ( .D(n392), .CK(clk), .Q(addrD[10]) );
  DFFHQ \driver/x_reg[0]  ( .D(n391), .CK(clk), .Q(addrD[6]) );
  DFFHQ \driver/x_reg[1]  ( .D(n390), .CK(clk), .Q(addrD[7]) );
  DFFHQ \driver/x_reg[2]  ( .D(n389), .CK(clk), .Q(addrD[8]) );
  DFFHQ \driver/x_reg[3]  ( .D(n388), .CK(clk), .Q(addrD[9]) );
  DFFHQ \driver/state_reg[0]  ( .D(n386), .CK(clk), .Q(state[0]) );
  EDFFTSHQ \driver/state_reg[1]  ( .SN(n367), .D(n448), .E(n729), .CK(clk), 
        .Q(state[1]) );
  DFFHQ \driver/state_reg[2]  ( .D(n387), .CK(clk), .Q(state[2]) );
  DFFHQ \driver/dori_o_reg  ( .D(n385), .CK(clk), .Q(dori_o) );
  DFFRHQ \decider/addrT_reg[0]  ( .D(n384), .CK(clk), .RN(rstn), .Q(addrT[0])
         );
  DFFRHQ \decider/addrT_reg[1]  ( .D(n383), .CK(clk), .RN(rstn), .Q(addrT[1])
         );
  DFFRHQ \decider/addrT_reg[2]  ( .D(n382), .CK(clk), .RN(rstn), .Q(addrT[2])
         );
  DFFRHQ \decider/addrT_reg[3]  ( .D(n381), .CK(clk), .RN(rstn), .Q(addrT[3])
         );
  DFFRHQ \decider/addrT_reg[4]  ( .D(n380), .CK(clk), .RN(rstn), .Q(addrT[4])
         );
  DFFRHQ \decider/addrT_reg[5]  ( .D(n379), .CK(clk), .RN(rstn), .Q(addrT[5])
         );
  DFFRHQ \decider/addrT_reg[6]  ( .D(n378), .CK(clk), .RN(rstn), .Q(addrT[6])
         );
  DFFRHQ \decider/addrT_reg[7]  ( .D(n377), .CK(clk), .RN(rstn), .Q(addrT[7])
         );
  DFFRHQ \decider/addrT_reg[8]  ( .D(n376), .CK(clk), .RN(rstn), .Q(addrT[8])
         );
  DFFRHQ \decider/addrT_reg[9]  ( .D(n375), .CK(clk), .RN(rstn), .Q(addrT[9])
         );
  DFFHQ \driver/db_o_reg[6]  ( .D(n368), .CK(clk), .Q(db_o[6]) );
  DFFHQ \driver/db_o_reg[5]  ( .D(n369), .CK(clk), .Q(db_o[5]) );
  DFFHQ \driver/db_o_reg[4]  ( .D(n370), .CK(clk), .Q(db_o[4]) );
  DFFHQ \driver/db_o_reg[3]  ( .D(n371), .CK(clk), .Q(db_o[3]) );
  DFFHQ \driver/db_o_reg[2]  ( .D(n372), .CK(clk), .Q(db_o[2]) );
  DFFHQ \driver/db_o_reg[1]  ( .D(n700), .CK(clk), .Q(db_o[1]) );
  DFFHQ \driver/db_o_reg[0]  ( .D(n701), .CK(clk), .Q(db_o[0]) );
  DFFHQ \driver/db_o_reg[7]  ( .D(n702), .CK(clk), .Q(db_o[7]) );
  DFFRHQ \clock_divider/cnt5k_reg[11]  ( .D(\clock_divider/N29 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[11] ) );
  DFFRHQ \clock_divider/cnt5k_reg[0]  ( .D(\clock_divider/N18 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[0] ) );
  DFFRHQ \clock_divider/cnt5k_reg[1]  ( .D(\clock_divider/N19 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[1] ) );
  DFFRHQ \clock_divider/cnt5k_reg[2]  ( .D(\clock_divider/N20 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[2] ) );
  DFFRHQ \clock_divider/cnt5k_reg[3]  ( .D(\clock_divider/N21 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[3] ) );
  DFFRHQ \clock_divider/cnt5k_reg[4]  ( .D(\clock_divider/N22 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[4] ) );
  DFFRHQ \clock_divider/cnt5k_reg[5]  ( .D(\clock_divider/N23 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[5] ) );
  DFFRHQ \clock_divider/cnt5k_reg[6]  ( .D(\clock_divider/N24 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[6] ) );
  DFFRHQ \clock_divider/cnt5k_reg[7]  ( .D(\clock_divider/N25 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[7] ) );
  DFFRHQ \clock_divider/cnt5k_reg[8]  ( .D(\clock_divider/N26 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[8] ) );
  DFFRHQ \clock_divider/cnt5k_reg[9]  ( .D(\clock_divider/N27 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[9] ) );
  DFFRHQ \clock_divider/cnt5k_reg[10]  ( .D(\clock_divider/N28 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[10] ) );
  OAI2BB2 U312 ( .B0(n452), .B1(n703), .A0N(\decider/N96 ), .A1N(n453), .Y(
        \U1/U2/Z_9 ) );
  OAI2BB2 U314 ( .B0(n454), .B1(n704), .A0N(\decider/N95 ), .A1N(n455), .Y(
        \U1/U2/Z_8 ) );
  OAI2BB2 U316 ( .B0(n452), .B1(n705), .A0N(\decider/N94 ), .A1N(n453), .Y(
        \U1/U2/Z_7 ) );
  OAI2BB2 U318 ( .B0(n454), .B1(n706), .A0N(\decider/N93 ), .A1N(n455), .Y(
        \U1/U2/Z_6 ) );
  OAI2BB2 U320 ( .B0(n452), .B1(n707), .A0N(\decider/N92 ), .A1N(n453), .Y(
        \U1/U2/Z_5 ) );
  OAI2BB2 U322 ( .B0(n454), .B1(n708), .A0N(\decider/N91 ), .A1N(n455), .Y(
        \U1/U2/Z_4 ) );
  OAI2BB2 U324 ( .B0(n452), .B1(n709), .A0N(\decider/N90 ), .A1N(n453), .Y(
        \U1/U2/Z_3 ) );
  OAI2BB2 U326 ( .B0(n454), .B1(n710), .A0N(\decider/N89 ), .A1N(n455), .Y(
        \U1/U2/Z_2 ) );
  OAI2BB2 U340 ( .B0(n452), .B1(n711), .A0N(\decider/N88 ), .A1N(n453), .Y(
        \U1/U2/Z_1 ) );
  OAI2BB2 U342 ( .B0(n454), .B1(n712), .A0N(\decider/N87 ), .A1N(n455), .Y(
        \U1/U2/Z_0 ) );
  ADDF \r250/U2_1  ( .A(\U1/U5/Z_1 ), .B(n727), .CI(\r250/carry[1] ), .CO(
        \r250/carry[2] ), .S(\decider/N88 ) );
  ADDF \r250/U2_2  ( .A(\U1/U5/Z_2 ), .B(n720), .CI(\r250/carry[2] ), .CO(
        \r250/carry[3] ), .S(\decider/N89 ) );
  ADDF \r250/U2_3  ( .A(\U1/U5/Z_3 ), .B(n719), .CI(\r250/carry[3] ), .CO(
        \r250/carry[4] ), .S(\decider/N90 ) );
  ADDF \r250/U2_4  ( .A(\U1/U5/Z_4 ), .B(n718), .CI(\r250/carry[4] ), .CO(
        \r250/carry[5] ), .S(\decider/N91 ) );
  ADDF \r250/U2_5  ( .A(\U1/U5/Z_5 ), .B(n717), .CI(\r250/carry[5] ), .CO(
        \r250/carry[6] ), .S(\decider/N92 ) );
  ADDF \r250/U2_6  ( .A(\U1/U5/Z_6 ), .B(n716), .CI(\r250/carry[6] ), .CO(
        \r250/carry[7] ), .S(\decider/N93 ) );
  ADDF \r250/U2_7  ( .A(\U1/U5/Z_7 ), .B(n715), .CI(\r250/carry[7] ), .CO(
        \r250/carry[8] ), .S(\decider/N94 ) );
  ADDF \r250/U2_8  ( .A(\U1/U5/Z_8 ), .B(n714), .CI(\r250/carry[8] ), .CO(
        \r250/carry[9] ), .S(\decider/N95 ) );
  ADDF \r250/U2_9  ( .A(\U1/U5/Z_9 ), .B(n713), .CI(\r250/carry[9] ), .CO(
        \r250/carry[10] ), .S(\decider/N96 ) );
  ADDF \r250/U2_10  ( .A(\U1/U5/Z_10 ), .B(n726), .CI(\r250/carry[10] ), .CO(
        \r250/carry[11] ), .S(\decider/N97 ) );
  ADDF \r250/U2_11  ( .A(\U1/U5/Z_11 ), .B(n725), .CI(\r250/carry[11] ), .CO(
        \r250/carry[12] ), .S(\decider/N98 ) );
  ADDF \r250/U2_12  ( .A(\U1/U5/Z_12 ), .B(n724), .CI(\r250/carry[12] ), .CO(
        \r250/carry[13] ), .S(\decider/N99 ) );
  ADDF \r250/U2_13  ( .A(\U1/U5/Z_13 ), .B(n723), .CI(\r250/carry[13] ), .CO(
        \r250/carry[14] ), .S(\decider/N100 ) );
  ADDF \r250/U2_14  ( .A(\U1/U5/Z_14 ), .B(n722), .CI(\r250/carry[14] ), .CO(
        \r250/carry[15] ), .S(\decider/N101 ) );
  ADDF \r250/U2_15  ( .A(\U1/U5/Z_15 ), .B(n721), .CI(\r250/carry[15] ), .S(
        \decider/N102 ) );
  ADDF \r191/U2_3  ( .A(addrD[6]), .B(\r191/B_not[3] ), .CI(\r191/carry[3] ), 
        .CO(\r191/carry[4] ), .S(\decider/obstacle_right [3]) );
  ADDF \r191/U2_4  ( .A(addrD[7]), .B(\r191/B_not[4] ), .CI(\r191/carry[4] ), 
        .CO(\r191/carry[5] ), .S(\decider/obstacle_right [4]) );
  ADDF \r191/U2_5  ( .A(addrD[8]), .B(\r191/B_not[5] ), .CI(\r191/carry[5] ), 
        .CO(\r191/carry[6] ), .S(\decider/obstacle_right [5]) );
  ADDF \r191/U2_6  ( .A(addrD[9]), .B(\r191/B_not[6] ), .CI(\r191/carry[6] ), 
        .CO(\r191/carry[7] ), .S(\decider/obstacle_right [6]) );
  ADDF \r191/U2_7  ( .A(addrD[10]), .B(\r191/B_not[7] ), .CI(\r191/carry[7] ), 
        .CO(\r191/carry[8] ), .S(\decider/obstacle_right [7]) );
  ADDF \r191/U2_8  ( .A(\driver/*Logic0* ), .B(\r191/B_not[8] ), .CI(
        \r191/carry[8] ), .CO(\r191/carry[9] ), .S(\decider/obstacle_right [8]) );
  ADDF \r191/U2_9  ( .A(\driver/*Logic0* ), .B(\r191/B_not[9] ), .CI(
        \r191/carry[9] ), .CO(\r191/carry[10] ), .S(
        \decider/obstacle_right [9]) );
  ADDF \r191/U2_10  ( .A(\driver/*Logic0* ), .B(\r191/B_not[10] ), .CI(
        \r191/carry[10] ), .CO(\r191/carry[11] ), .S(
        \decider/obstacle_right [10]) );
  ADDF \r191/U2_11  ( .A(\driver/*Logic0* ), .B(\r191/B_not[11] ), .CI(
        \r191/carry[11] ), .CO(\r191/carry[12] ), .S(
        \decider/obstacle_right [11]) );
  ADDF \r191/U2_12  ( .A(\driver/*Logic0* ), .B(\r191/B_not[12] ), .CI(
        \r191/carry[12] ), .CO(\r191/carry[13] ), .S(
        \decider/obstacle_right [12]) );
  ADDF \r191/U2_13  ( .A(\driver/*Logic0* ), .B(\r191/B_not[13] ), .CI(
        \r191/carry[13] ), .CO(\r191/carry[14] ), .S(
        \decider/obstacle_right [13]) );
  ADDF \r191/U2_14  ( .A(\driver/*Logic0* ), .B(\r191/B_not[14] ), .CI(
        \r191/carry[14] ), .CO(\r191/carry[15] ), .S(
        \decider/obstacle_right [14]) );
  ADDF \r191/U2_15  ( .A(\driver/*Logic0* ), .B(\r191/B_not[15] ), .CI(
        \r191/carry[15] ), .S(\decider/obstacle_right [15]) );
  ADDF \r187/U2_0  ( .A(n731), .B(\r187/B_not[0] ), .CI(n736), .CO(
        \r187/carry[1] ), .S(\decider/rex_top [0]) );
  ADDF \r187/U2_1  ( .A(n732), .B(\r187/B_not[1] ), .CI(\r187/carry[1] ), .CO(
        \r187/carry[2] ), .S(\decider/rex_top [1]) );
  ADDF \r187/U2_2  ( .A(n733), .B(\r187/B_not[2] ), .CI(\r187/carry[2] ), .CO(
        \r187/carry[3] ), .S(\decider/rex_top [2]) );
  ADDF \r187/U2_3  ( .A(n734), .B(\r187/B_not[3] ), .CI(\r187/carry[3] ), .CO(
        \r187/carry[4] ), .S(\decider/rex_top [3]) );
  ADDF \r187/U2_4  ( .A(n735), .B(\r187/B_not[4] ), .CI(\r187/carry[4] ), .CO(
        \r187/carry[5] ), .S(\decider/rex_top [4]) );
  ADDF \r187/U2_5  ( .A(n730), .B(\r187/B_not[5] ), .CI(\r187/carry[5] ), .CO(
        \r187/carry[6] ), .S(\decider/rex_top [5]) );
  ADDF \r187/U2_6  ( .A(\driver/*Logic0* ), .B(\r187/B_not[6] ), .CI(
        \r187/carry[6] ), .CO(\r187/carry[7] ), .S(\decider/rex_top [6]) );
  ADDF \r187/U2_7  ( .A(\driver/*Logic0* ), .B(\r187/B_not[7] ), .CI(
        \r187/carry[7] ), .CO(\r187/carry[8] ), .S(\decider/rex_top [7]) );
  ADDF \r187/U2_8  ( .A(\driver/*Logic0* ), .B(\r187/B_not[8] ), .CI(
        \r187/carry[8] ), .CO(\r187/carry[9] ), .S(\decider/rex_top [8]) );
  ADDF \r187/U2_9  ( .A(\driver/*Logic0* ), .B(\r187/B_not[9] ), .CI(
        \r187/carry[9] ), .CO(\r187/carry[10] ), .S(\decider/rex_top [9]) );
  ADDF \r187/U2_10  ( .A(\driver/*Logic0* ), .B(\r187/B_not[10] ), .CI(
        \r187/carry[10] ), .CO(\r187/carry[11] ), .S(\decider/rex_top [10]) );
  ADDF \r187/U2_11  ( .A(\driver/*Logic0* ), .B(\r187/B_not[11] ), .CI(
        \r187/carry[11] ), .CO(\r187/carry[12] ), .S(\decider/rex_top [11]) );
  ADDF \r187/U2_12  ( .A(\driver/*Logic0* ), .B(\r187/B_not[12] ), .CI(
        \r187/carry[12] ), .CO(\r187/carry[13] ), .S(\decider/rex_top [12]) );
  ADDF \r187/U2_13  ( .A(\driver/*Logic0* ), .B(\r187/B_not[13] ), .CI(
        \r187/carry[13] ), .CO(\r187/carry[14] ), .S(\decider/rex_top [13]) );
  ADDF \r187/U2_14  ( .A(\driver/*Logic0* ), .B(\r187/B_not[14] ), .CI(
        \r187/carry[14] ), .CO(\r187/carry[15] ), .S(\decider/rex_top [14]) );
  ADDF \r187/U2_15  ( .A(\driver/*Logic0* ), .B(\r187/B_not[15] ), .CI(
        \r187/carry[15] ), .S(\decider/rex_top [15]) );
  ADDF \r62/S3_2_3  ( .A(\U1/U3/Z_2 ), .B(n444), .CI(\U1/U3/Z_1 ), .CO(
        \r62/CARRYB[2][3] ), .S(\r62/SUMB[2][3] ) );
  ADDF \r62/S2_2_2  ( .A(\r62/ab[2][2] ), .B(n443), .CI(\r62/SUMB[1][3] ), 
        .CO(\r62/CARRYB[2][2] ), .S(\r62/SUMB[2][2] ) );
  ADDF \r62/S3_3_3  ( .A(\U1/U3/Z_3 ), .B(\r62/CARRYB[2][3] ), .CI(\U1/U3/Z_2 ), .CO(\r62/CARRYB[3][3] ), .S(\r62/SUMB[3][3] ) );
  ADDF \r62/S2_3_2  ( .A(\r62/ab[3][2] ), .B(\r62/CARRYB[2][2] ), .CI(
        \r62/SUMB[2][3] ), .CO(\r62/CARRYB[3][2] ), .S(\r62/SUMB[3][2] ) );
  ADDF \r62/S1_3_0  ( .A(\r62/ab[3][0] ), .B(n442), .CI(\r62/SUMB[1][2] ), 
        .CO(\r62/CARRYB[3][0] ), .S(\decider/N58 ) );
  ADDF \r62/S3_4_3  ( .A(\U1/U3/Z_4 ), .B(\r62/CARRYB[3][3] ), .CI(\U1/U3/Z_3 ), .CO(\r62/CARRYB[4][3] ), .S(\r62/SUMB[4][3] ) );
  ADDF \r62/S2_4_2  ( .A(\r62/ab[4][2] ), .B(\r62/CARRYB[3][2] ), .CI(
        \r62/SUMB[3][3] ), .CO(\r62/CARRYB[4][2] ), .S(\r62/SUMB[4][2] ) );
  ADDF \r62/S1_4_0  ( .A(\r62/ab[4][0] ), .B(\r62/CARRYB[3][0] ), .CI(
        \r62/SUMB[2][2] ), .CO(\r62/CARRYB[4][0] ), .S(\r62/PROD1[4] ) );
  ADDF \r62/S3_5_3  ( .A(\r62/ab[5][2] ), .B(\r62/CARRYB[4][3] ), .CI(
        \U1/U3/Z_4 ), .CO(\r62/CARRYB[5][3] ), .S(\r62/SUMB[5][3] ) );
  ADDF \r62/S2_5_2  ( .A(\r62/ab[5][2] ), .B(\r62/CARRYB[4][2] ), .CI(
        \r62/SUMB[4][3] ), .CO(\r62/CARRYB[5][2] ), .S(\r62/SUMB[5][2] ) );
  ADDF \r62/S3_6_3  ( .A(\r62/ab[6][2] ), .B(\r62/CARRYB[5][3] ), .CI(
        \r62/ab[5][2] ), .CO(\r62/CARRYB[6][3] ), .S(\r62/SUMB[6][3] ) );
  ADDF \r62/S2_6_2  ( .A(\r62/ab[6][2] ), .B(\r62/CARRYB[5][2] ), .CI(
        \r62/SUMB[5][3] ), .CO(\r62/CARRYB[6][2] ), .S(\r62/SUMB[6][2] ) );
  ADDF \r62/S3_7_3  ( .A(\r62/ab[7][2] ), .B(\r62/CARRYB[6][3] ), .CI(
        \r62/ab[6][2] ), .CO(\r62/CARRYB[7][3] ), .S(\r62/SUMB[7][3] ) );
  ADDF \r62/S2_7_2  ( .A(\r62/ab[7][2] ), .B(\r62/CARRYB[6][2] ), .CI(
        \r62/SUMB[6][3] ), .CO(\r62/CARRYB[7][2] ), .S(\r62/SUMB[7][2] ) );
  ADDF \r62/S3_8_3  ( .A(\r62/ab[8][2] ), .B(\r62/CARRYB[7][3] ), .CI(
        \r62/ab[7][2] ), .CO(\r62/CARRYB[8][3] ), .S(\r62/SUMB[8][3] ) );
  ADDF \r62/S2_8_2  ( .A(\r62/ab[8][2] ), .B(\r62/CARRYB[7][2] ), .CI(
        \r62/SUMB[7][3] ), .CO(\r62/CARRYB[8][2] ), .S(\r62/SUMB[8][2] ) );
  ADDF \r62/S3_9_3  ( .A(\r62/ab[9][2] ), .B(\r62/CARRYB[8][3] ), .CI(
        \r62/ab[8][2] ), .CO(\r62/CARRYB[9][3] ), .S(\r62/SUMB[9][3] ) );
  ADDF \r62/S2_9_2  ( .A(\r62/ab[9][2] ), .B(\r62/CARRYB[8][2] ), .CI(
        \r62/SUMB[8][3] ), .CO(\r62/CARRYB[9][2] ), .S(\r62/SUMB[9][2] ) );
  ADDF \r62/S3_10_3  ( .A(\r62/ab[10][2] ), .B(\r62/CARRYB[9][3] ), .CI(
        \r62/ab[9][2] ), .CO(\r62/CARRYB[10][3] ), .S(\r62/SUMB[10][3] ) );
  ADDF \r62/S2_10_2  ( .A(\r62/ab[10][2] ), .B(\r62/CARRYB[9][2] ), .CI(
        \r62/SUMB[9][3] ), .CO(\r62/CARRYB[10][2] ), .S(\r62/SUMB[10][2] ) );
  ADDF \r62/S3_11_3  ( .A(\r62/ab[11][2] ), .B(\r62/CARRYB[10][3] ), .CI(
        \r62/ab[10][2] ), .CO(\r62/CARRYB[11][3] ), .S(\r62/SUMB[11][3] ) );
  ADDF \r62/S2_11_2  ( .A(\r62/ab[11][2] ), .B(\r62/CARRYB[10][2] ), .CI(
        \r62/SUMB[10][3] ), .CO(\r62/CARRYB[11][2] ), .S(\r62/SUMB[11][2] ) );
  ADDF \r62/S5_3  ( .A(\r62/ab[12][2] ), .B(\r62/CARRYB[11][3] ), .CI(
        \r62/ab[11][2] ), .S(\r62/SUMB[12][3] ) );
  ADDF \r62/S4_2  ( .A(\r62/ab[12][2] ), .B(\r62/CARRYB[11][2] ), .CI(
        \r62/SUMB[11][3] ), .CO(\r62/CARRYB[12][2] ), .S(\r62/SUMB[12][2] ) );
  ADDF \r50/U1_1  ( .A(n406), .B(\U1/U2/Z_1 ), .CI(n441), .CO(\r50/carry[2] ), 
        .S(\decider/N85 ) );
  ADDF \r50/U1_3  ( .A(n406), .B(\U1/U2/Z_3 ), .CI(n440), .CO(\r50/carry[4] ), 
        .S(\decider/N83 ) );
  ADDF \r50/U1_6  ( .A(n406), .B(\U1/U2/Z_6 ), .CI(n439), .CO(\r50/carry[7] ), 
        .S(\decider/N80 ) );
  AND2 U345 ( .A(\decider/rex_top [3]), .B(
        \sub_0_root_decider/sub_49/carry[3] ), .Y(n402) );
  AND2 U346 ( .A(\r62/SUMB[10][2] ), .B(n430), .Y(n403) );
  AND2 U347 ( .A(n434), .B(\r62/SUMB[7][2] ), .Y(n404) );
  OR2 U348 ( .A(n455), .B(n457), .Y(n405) );
  NAND4 U349 ( .A(cs_o[0]), .B(n699), .C(\decider/sub_45/carry[5] ), .D(
        \decider/posy_m_rex_top[15] ), .Y(n406) );
  AND2 U350 ( .A(n734), .B(n733), .Y(n407) );
  AND2 U351 ( .A(\clock_divider/cnt5k[1] ), .B(\clock_divider/cnt5k[0] ), .Y(
        n408) );
  AND2 U352 ( .A(\clock_divider/cnt5k[2] ), .B(n408), .Y(n409) );
  AND2 U353 ( .A(\clock_divider/cnt5k[3] ), .B(n409), .Y(n410) );
  AND2 U354 ( .A(\clock_divider/cnt5k[4] ), .B(n410), .Y(n411) );
  AND2 U355 ( .A(\clock_divider/cnt5k[5] ), .B(n411), .Y(n412) );
  AND2 U356 ( .A(\clock_divider/cnt5k[6] ), .B(n412), .Y(n413) );
  AND2 U357 ( .A(\clock_divider/cnt5k[7] ), .B(n413), .Y(n414) );
  AND2 U358 ( .A(\clock_divider/cnt5k[8] ), .B(n414), .Y(n415) );
  AND2 U359 ( .A(\clock_divider/cnt5k[9] ), .B(n415), .Y(n416) );
  AND2 U360 ( .A(\clock_divider/cnt5k[10] ), .B(n416), .Y(n417) );
  AND2 U361 ( .A(addrD[7]), .B(addrD[6]), .Y(n418) );
  AND2 U362 ( .A(addrD[8]), .B(n418), .Y(n419) );
  AND2 U363 ( .A(\U1/U2/Z_4 ), .B(\r50/carry[4] ), .Y(n420) );
  AND2 U364 ( .A(\U1/U2/Z_7 ), .B(\r50/carry[7] ), .Y(n421) );
  AND2 U365 ( .A(\U1/U2/Z_8 ), .B(n421), .Y(n422) );
  AND2 U366 ( .A(\U1/U2/Z_9 ), .B(n422), .Y(n423) );
  AND2 U367 ( .A(\U1/U2/Z_10 ), .B(n423), .Y(n424) );
  AND2 U368 ( .A(\U1/U2/Z_11 ), .B(n424), .Y(n425) );
  AND2 U369 ( .A(\U1/U2/Z_12 ), .B(n425), .Y(n426) );
  AND2 U370 ( .A(\U1/U2/Z_13 ), .B(n426), .Y(n427) );
  AND2 U371 ( .A(n403), .B(\r62/SUMB[11][2] ), .Y(n428) );
  AND2 U372 ( .A(n404), .B(\r62/SUMB[8][2] ), .Y(n429) );
  AND2 U373 ( .A(n429), .B(\r62/SUMB[9][2] ), .Y(n430) );
  AND2 U374 ( .A(\r62/CARRYB[4][0] ), .B(\r62/SUMB[3][2] ), .Y(n431) );
  AND2 U375 ( .A(n431), .B(\r62/SUMB[4][2] ), .Y(n432) );
  AND2 U376 ( .A(n432), .B(\r62/SUMB[5][2] ), .Y(n433) );
  AND2 U377 ( .A(n433), .B(\r62/SUMB[6][2] ), .Y(n434) );
  XOR2 U378 ( .A(\decider/obstacle_right [15]), .B(
        \sub_0_root_decider/sub_73/carry[15] ), .Y(n435) );
  AND2 U379 ( .A(\clock_divider/cnt5k[11] ), .B(n417), .Y(n436) );
  AND2 U380 ( .A(addrD[9]), .B(n419), .Y(n437) );
  AND2 U381 ( .A(\U1/U2/Z_14 ), .B(n427), .Y(n438) );
  AND2 U382 ( .A(\U1/U2/Z_5 ), .B(n420), .Y(n439) );
  AND2 U383 ( .A(\U1/U2/Z_2 ), .B(\r50/carry[2] ), .Y(n440) );
  AND2 U384 ( .A(\U1/U2/Z_0 ), .B(n406), .Y(n441) );
  AND2 U385 ( .A(\r62/ab[2][0] ), .B(\r62/ab[0][2] ), .Y(n442) );
  AND2 U386 ( .A(\U1/U3/Z_0 ), .B(\r62/ab[1][2] ), .Y(n443) );
  AND2 U387 ( .A(\U1/U3/Z_0 ), .B(\U1/U3/Z_1 ), .Y(n444) );
  INV U388 ( .A(n586), .Y(n445) );
  INV U389 ( .A(n445), .Y(n446) );
  INV U390 ( .A(n366), .Y(n447) );
  INV U391 ( .A(n447), .Y(n448) );
  INV U392 ( .A(n405), .Y(n449) );
  INV U393 ( .A(n559), .Y(n450) );
  INV U394 ( .A(n450), .Y(n451) );
  INV U395 ( .A(n406), .Y(n452) );
  INV U396 ( .A(n406), .Y(n453) );
  INV U397 ( .A(n406), .Y(n454) );
  INV U398 ( .A(n406), .Y(n455) );
  INV U399 ( .A(n604), .Y(n456) );
  INV U400 ( .A(n456), .Y(n457) );
  BUF U401 ( .I(n498), .O(n458) );
  LOGIC_0 U402 ( .LOGIC_0_PIN(\driver/*Logic0* ) );
  LOGIC_1 U403 ( .LOGIC_1_PIN(n736) );
  NAND2 U404 ( .A(addrD[5]), .B(n488), .Y(\decider/sub_75/carry[6] ) );
  XNOR2 U405 ( .A(n730), .B(\decider/sub_75/carry[5] ), .Y(
        \decider/posy_m_obstacle_top [5]) );
  NAND2 U406 ( .A(n459), .B(n460), .Y(\sub_0_root_decider/sub_49/carry[11] )
         );
  XNOR2 U407 ( .A(\decider/rex_top [10]), .B(
        \sub_0_root_decider/sub_49/carry[10] ), .Y(
        \decider/posy_m_rex_top[10] ) );
  INV U408 ( .A(\decider/rex_top [10]), .Y(n459) );
  INV U409 ( .A(\sub_0_root_decider/sub_49/carry[10] ), .Y(n460) );
  NAND2 U410 ( .A(n461), .B(n462), .Y(\sub_0_root_decider/sub_49/carry[12] )
         );
  XNOR2 U411 ( .A(\decider/rex_top [11]), .B(
        \sub_0_root_decider/sub_49/carry[11] ), .Y(
        \decider/posy_m_rex_top[11] ) );
  INV U412 ( .A(\decider/rex_top [11]), .Y(n461) );
  INV U413 ( .A(\sub_0_root_decider/sub_49/carry[11] ), .Y(n462) );
  NAND2 U414 ( .A(n463), .B(n464), .Y(\sub_0_root_decider/sub_49/carry[13] )
         );
  XNOR2 U415 ( .A(\decider/rex_top [12]), .B(
        \sub_0_root_decider/sub_49/carry[12] ), .Y(
        \decider/posy_m_rex_top[12] ) );
  INV U416 ( .A(\decider/rex_top [12]), .Y(n463) );
  INV U417 ( .A(\sub_0_root_decider/sub_49/carry[12] ), .Y(n464) );
  NAND2 U418 ( .A(n465), .B(n466), .Y(\sub_0_root_decider/sub_49/carry[14] )
         );
  XNOR2 U419 ( .A(\decider/rex_top [13]), .B(
        \sub_0_root_decider/sub_49/carry[13] ), .Y(
        \decider/posy_m_rex_top[13] ) );
  INV U420 ( .A(\decider/rex_top [13]), .Y(n465) );
  INV U421 ( .A(\sub_0_root_decider/sub_49/carry[13] ), .Y(n466) );
  NAND2 U422 ( .A(n467), .B(n468), .Y(\sub_0_root_decider/sub_49/carry[15] )
         );
  XNOR2 U423 ( .A(\decider/rex_top [14]), .B(
        \sub_0_root_decider/sub_49/carry[14] ), .Y(
        \decider/posy_m_rex_top[14] ) );
  INV U424 ( .A(\decider/rex_top [14]), .Y(n467) );
  INV U425 ( .A(\sub_0_root_decider/sub_49/carry[14] ), .Y(n468) );
  XNOR2 U426 ( .A(\decider/rex_top [15]), .B(
        \sub_0_root_decider/sub_49/carry[15] ), .Y(
        \decider/posy_m_rex_top[15] ) );
  NAND2 U427 ( .A(n469), .B(n470), .Y(\sub_0_root_decider/sub_49/carry[2] ) );
  XNOR2 U428 ( .A(\decider/rex_top [1]), .B(\decider/rex_top [0]), .Y(
        \decider/posy_m_rex_top[1] ) );
  INV U429 ( .A(\decider/rex_top [1]), .Y(n469) );
  INV U430 ( .A(\decider/rex_top [0]), .Y(n470) );
  NAND2 U431 ( .A(n471), .B(n472), .Y(\sub_0_root_decider/sub_49/carry[3] ) );
  XNOR2 U432 ( .A(\decider/rex_top [2]), .B(
        \sub_0_root_decider/sub_49/carry[2] ), .Y(\decider/posy_m_rex_top[2] )
         );
  INV U433 ( .A(\decider/rex_top [2]), .Y(n471) );
  INV U434 ( .A(\sub_0_root_decider/sub_49/carry[2] ), .Y(n472) );
  NAND2 U435 ( .A(n473), .B(n489), .Y(\sub_0_root_decider/sub_49/carry[6] ) );
  XNOR2 U436 ( .A(\decider/rex_top [5]), .B(
        \sub_0_root_decider/sub_49/carry[5] ), .Y(\decider/posy_m_rex_top[5] )
         );
  INV U437 ( .A(\decider/rex_top [5]), .Y(n473) );
  NAND2 U438 ( .A(n474), .B(n475), .Y(\sub_0_root_decider/sub_49/carry[7] ) );
  XNOR2 U439 ( .A(\decider/rex_top [6]), .B(
        \sub_0_root_decider/sub_49/carry[6] ), .Y(\decider/posy_m_rex_top[6] )
         );
  INV U440 ( .A(\decider/rex_top [6]), .Y(n474) );
  INV U441 ( .A(\sub_0_root_decider/sub_49/carry[6] ), .Y(n475) );
  NAND2 U442 ( .A(n476), .B(n477), .Y(\sub_0_root_decider/sub_49/carry[8] ) );
  XNOR2 U443 ( .A(\decider/rex_top [7]), .B(
        \sub_0_root_decider/sub_49/carry[7] ), .Y(\decider/posy_m_rex_top[7] )
         );
  INV U444 ( .A(\decider/rex_top [7]), .Y(n476) );
  INV U445 ( .A(\sub_0_root_decider/sub_49/carry[7] ), .Y(n477) );
  NAND2 U446 ( .A(n478), .B(n479), .Y(\sub_0_root_decider/sub_49/carry[9] ) );
  XNOR2 U447 ( .A(\decider/rex_top [8]), .B(
        \sub_0_root_decider/sub_49/carry[8] ), .Y(\decider/posy_m_rex_top[8] )
         );
  INV U448 ( .A(\decider/rex_top [8]), .Y(n478) );
  INV U449 ( .A(\sub_0_root_decider/sub_49/carry[8] ), .Y(n479) );
  NAND2 U450 ( .A(n480), .B(n481), .Y(\sub_0_root_decider/sub_49/carry[10] )
         );
  XNOR2 U451 ( .A(\decider/rex_top [9]), .B(
        \sub_0_root_decider/sub_49/carry[9] ), .Y(\decider/posy_m_rex_top[9] )
         );
  INV U452 ( .A(\decider/rex_top [9]), .Y(n480) );
  INV U453 ( .A(\sub_0_root_decider/sub_49/carry[9] ), .Y(n481) );
  NAND2 U454 ( .A(n482), .B(n483), .Y(\r250/carry[1] ) );
  XNOR2 U455 ( .A(n728), .B(\U1/U5/Z_0 ), .Y(\decider/N87 ) );
  INV U456 ( .A(n728), .Y(n482) );
  INV U457 ( .A(\U1/U5/Z_0 ), .Y(n483) );
  NAND2 U458 ( .A(n585), .B(n484), .Y(\decider/sub_45/carry[5] ) );
  XNOR2 U459 ( .A(addrD[10]), .B(\decider/sub_45/carry[4] ), .Y(
        \decider/posx_m_rex_left [7]) );
  INV U460 ( .A(\decider/sub_45/carry[4] ), .Y(n484) );
  NAND2 U461 ( .A(n590), .B(n485), .Y(\decider/sub_45/carry[4] ) );
  XNOR2 U462 ( .A(addrD[9]), .B(\decider/sub_45/carry[3] ), .Y(
        \decider/posx_m_rex_left [6]) );
  INV U463 ( .A(\decider/sub_45/carry[3] ), .Y(n485) );
  NAND2 U464 ( .A(n589), .B(n486), .Y(\decider/sub_45/carry[3] ) );
  XNOR2 U465 ( .A(addrD[8]), .B(\decider/sub_45/carry[2] ), .Y(
        \decider/posx_m_rex_left [5]) );
  INV U466 ( .A(\decider/sub_45/carry[2] ), .Y(n486) );
  NAND2 U467 ( .A(n588), .B(n487), .Y(\decider/sub_45/carry[2] ) );
  XNOR2 U468 ( .A(addrD[7]), .B(addrD[6]), .Y(\decider/posx_m_rex_left [4]) );
  INV U469 ( .A(addrD[6]), .Y(n487) );
  XOR2 U470 ( .A(n734), .B(n733), .Y(\decider/posy_m_obstacle_top [3]) );
  XOR2 U471 ( .A(n735), .B(n407), .Y(\decider/posy_m_obstacle_top [4]) );
  NAND2 U472 ( .A(n735), .B(n407), .Y(n488) );
  INV U473 ( .A(n488), .Y(\decider/sub_75/carry[5] ) );
  XOR2 U474 ( .A(\clock_divider/cnt5k[1] ), .B(\clock_divider/cnt5k[0] ), .Y(
        \clock_divider/N6 ) );
  XOR2 U475 ( .A(\clock_divider/cnt5k[2] ), .B(n408), .Y(\clock_divider/N7 )
         );
  XOR2 U476 ( .A(\clock_divider/cnt5k[3] ), .B(n409), .Y(\clock_divider/N8 )
         );
  XOR2 U477 ( .A(\clock_divider/cnt5k[4] ), .B(n410), .Y(\clock_divider/N9 )
         );
  XOR2 U478 ( .A(\clock_divider/cnt5k[5] ), .B(n411), .Y(\clock_divider/N10 )
         );
  XOR2 U479 ( .A(\clock_divider/cnt5k[6] ), .B(n412), .Y(\clock_divider/N11 )
         );
  XOR2 U480 ( .A(\clock_divider/cnt5k[7] ), .B(n413), .Y(\clock_divider/N12 )
         );
  XOR2 U481 ( .A(\clock_divider/cnt5k[8] ), .B(n414), .Y(\clock_divider/N13 )
         );
  XOR2 U482 ( .A(\clock_divider/cnt5k[9] ), .B(n415), .Y(\clock_divider/N14 )
         );
  XOR2 U483 ( .A(\clock_divider/cnt5k[10] ), .B(n416), .Y(\clock_divider/N15 )
         );
  XOR2 U484 ( .A(\clock_divider/cnt5k[11] ), .B(n417), .Y(\clock_divider/N16 )
         );
  XOR2 U485 ( .A(\clock_divider/cnt5k[12] ), .B(n436), .Y(\clock_divider/N17 )
         );
  XOR2 U486 ( .A(addrD[7]), .B(addrD[6]), .Y(\driver/N44 ) );
  XOR2 U487 ( .A(addrD[8]), .B(n418), .Y(\driver/N45 ) );
  XOR2 U488 ( .A(addrD[9]), .B(n419), .Y(\driver/N46 ) );
  XOR2 U489 ( .A(addrD[10]), .B(n437), .Y(\driver/N47 ) );
  XOR2 U490 ( .A(\decider/rex_top [3]), .B(
        \sub_0_root_decider/sub_49/carry[3] ), .Y(\decider/posy_m_rex_top[3] )
         );
  XOR2 U491 ( .A(\decider/rex_top [4]), .B(n402), .Y(
        \decider/posy_m_rex_top[4] ) );
  NAND2 U492 ( .A(\decider/rex_top [4]), .B(n402), .Y(n489) );
  INV U493 ( .A(n489), .Y(\sub_0_root_decider/sub_49/carry[5] ) );
  XOR2 U494 ( .A(n403), .B(\r62/SUMB[11][2] ), .Y(\r62/A1[11] ) );
  XOR2 U495 ( .A(\r62/CARRYB[12][2] ), .B(\r62/SUMB[12][3] ), .Y(\r62/A1[13] )
         );
  XOR2 U496 ( .A(\r62/ab[1][2] ), .B(\U1/U3/Z_0 ), .Y(\r62/SUMB[1][2] ) );
  XOR2 U497 ( .A(\U1/U3/Z_1 ), .B(\U1/U3/Z_0 ), .Y(\r62/SUMB[1][3] ) );
  XOR2 U498 ( .A(\U1/U2/Z_0 ), .B(n406), .Y(\decider/N86 ) );
  XOR2 U499 ( .A(\U1/U2/Z_2 ), .B(\r50/carry[2] ), .Y(\decider/N84 ) );
  XOR2 U500 ( .A(\U1/U2/Z_4 ), .B(\r50/carry[4] ), .Y(\decider/N82 ) );
  XOR2 U501 ( .A(\U1/U2/Z_5 ), .B(n420), .Y(\decider/N81 ) );
  XOR2 U502 ( .A(\U1/U2/Z_7 ), .B(\r50/carry[7] ), .Y(\decider/N79 ) );
  XOR2 U503 ( .A(\U1/U2/Z_8 ), .B(n421), .Y(\decider/N78 ) );
  XOR2 U504 ( .A(\U1/U2/Z_9 ), .B(n422), .Y(\decider/N77 ) );
  XOR2 U505 ( .A(\U1/U2/Z_10 ), .B(n423), .Y(\decider/N76 ) );
  XOR2 U506 ( .A(\U1/U2/Z_11 ), .B(n424), .Y(\decider/N75 ) );
  XOR2 U507 ( .A(\U1/U2/Z_12 ), .B(n425), .Y(\decider/N74 ) );
  XOR2 U508 ( .A(\U1/U2/Z_13 ), .B(n426), .Y(\decider/N73 ) );
  XOR2 U509 ( .A(\U1/U2/Z_14 ), .B(n427), .Y(\decider/N72 ) );
  XOR2 U510 ( .A(\U1/U2/Z_15 ), .B(n438), .Y(\decider/N71 ) );
  XOR2 U511 ( .A(\r62/ab[2][0] ), .B(\r62/ab[0][2] ), .Y(\decider/N57 ) );
  XOR2 U512 ( .A(n404), .B(\r62/SUMB[8][2] ), .Y(\decider/N65 ) );
  XOR2 U513 ( .A(n429), .B(\r62/SUMB[9][2] ), .Y(\r62/A1[9] ) );
  XOR2 U514 ( .A(n430), .B(\r62/SUMB[10][2] ), .Y(\r62/SUMB[12][0] ) );
  XOR2 U515 ( .A(\r62/CARRYB[4][0] ), .B(\r62/SUMB[3][2] ), .Y(\decider/N60 )
         );
  XOR2 U516 ( .A(n431), .B(\r62/SUMB[4][2] ), .Y(\decider/N61 ) );
  XOR2 U517 ( .A(n432), .B(\r62/SUMB[5][2] ), .Y(\decider/N62 ) );
  XOR2 U518 ( .A(n433), .B(\r62/SUMB[6][2] ), .Y(\decider/N63 ) );
  XOR2 U519 ( .A(n434), .B(\r62/SUMB[7][2] ), .Y(\decider/N64 ) );
  NAND2 U520 ( .A(n490), .B(n491), .Y(\sub_0_root_decider/sub_73/carry[15] )
         );
  NOR4B U521 ( .AN(n492), .B(\decider/obstacle_right [6]), .C(
        \decider/obstacle_right [4]), .D(\decider/obstacle_right [5]), .Y(n491) );
  NOR3 U522 ( .A(\decider/obstacle_right [7]), .B(\decider/obstacle_right [9]), 
        .C(\decider/obstacle_right [8]), .Y(n492) );
  NOR4B U523 ( .AN(n493), .B(\decider/obstacle_right [12]), .C(
        \decider/obstacle_right [11]), .D(\decider/obstacle_right [10]), .Y(
        n490) );
  NOR2 U524 ( .A(\decider/obstacle_right [14]), .B(
        \decider/obstacle_right [13]), .Y(n493) );
  NOR2B U525 ( .AN(\U1/U3/Z_4 ), .B(n454), .Y(\r62/ab[4][2] ) );
  NOR2B U526 ( .AN(\U1/U3/Z_4 ), .B(n406), .Y(\r62/ab[4][0] ) );
  NOR2B U527 ( .AN(\U1/U3/Z_3 ), .B(n455), .Y(\r62/ab[3][2] ) );
  NOR2B U528 ( .AN(\U1/U3/Z_3 ), .B(n406), .Y(\r62/ab[3][0] ) );
  NOR2B U529 ( .AN(\U1/U3/Z_2 ), .B(n452), .Y(\r62/ab[2][2] ) );
  NOR2B U530 ( .AN(\U1/U3/Z_2 ), .B(n406), .Y(\r62/ab[2][0] ) );
  NOR2B U531 ( .AN(\U1/U3/Z_1 ), .B(n453), .Y(\r62/ab[1][2] ) );
  NOR2B U532 ( .AN(\U1/U3/Z_0 ), .B(n454), .Y(\r62/ab[0][2] ) );
  NOR3 U533 ( .A(obstacle_left[0]), .B(obstacle_left[2]), .C(obstacle_left[1]), 
        .Y(\r191/carry[3] ) );
  INV U534 ( .A(obstacle_left[9]), .Y(\r191/B_not[9] ) );
  INV U535 ( .A(obstacle_left[8]), .Y(\r191/B_not[8] ) );
  INV U536 ( .A(obstacle_left[7]), .Y(\r191/B_not[7] ) );
  INV U537 ( .A(obstacle_left[6]), .Y(\r191/B_not[6] ) );
  INV U538 ( .A(obstacle_left[5]), .Y(\r191/B_not[5] ) );
  INV U539 ( .A(obstacle_left[4]), .Y(\r191/B_not[4] ) );
  INV U540 ( .A(obstacle_left[3]), .Y(\r191/B_not[3] ) );
  INV U541 ( .A(obstacle_left[15]), .Y(\r191/B_not[15] ) );
  INV U542 ( .A(obstacle_left[14]), .Y(\r191/B_not[14] ) );
  INV U543 ( .A(obstacle_left[13]), .Y(\r191/B_not[13] ) );
  INV U544 ( .A(obstacle_left[12]), .Y(\r191/B_not[12] ) );
  INV U545 ( .A(obstacle_left[11]), .Y(\r191/B_not[11] ) );
  INV U546 ( .A(obstacle_left[10]), .Y(\r191/B_not[10] ) );
  INV U547 ( .A(rex_down[9]), .Y(\r187/B_not[9] ) );
  INV U548 ( .A(rex_down[8]), .Y(\r187/B_not[8] ) );
  INV U549 ( .A(rex_down[7]), .Y(\r187/B_not[7] ) );
  INV U550 ( .A(rex_down[6]), .Y(\r187/B_not[6] ) );
  INV U551 ( .A(rex_down[5]), .Y(\r187/B_not[5] ) );
  INV U552 ( .A(rex_down[4]), .Y(\r187/B_not[4] ) );
  INV U553 ( .A(rex_down[3]), .Y(\r187/B_not[3] ) );
  INV U554 ( .A(rex_down[2]), .Y(\r187/B_not[2] ) );
  INV U555 ( .A(rex_down[1]), .Y(\r187/B_not[1] ) );
  INV U556 ( .A(rex_down[15]), .Y(\r187/B_not[15] ) );
  INV U557 ( .A(rex_down[14]), .Y(\r187/B_not[14] ) );
  INV U558 ( .A(rex_down[13]), .Y(\r187/B_not[13] ) );
  INV U559 ( .A(rex_down[12]), .Y(\r187/B_not[12] ) );
  INV U560 ( .A(rex_down[11]), .Y(\r187/B_not[11] ) );
  INV U561 ( .A(rex_down[10]), .Y(\r187/B_not[10] ) );
  INV U562 ( .A(rex_down[0]), .Y(\r187/B_not[0] ) );
  OAI211 U563 ( .A0(n494), .A1(n495), .B0(n496), .C0(n497), .Y(n700) );
  AOI222 U564 ( .A0(db_o[1]), .A1(n458), .B0(addrD[7]), .B1(n499), .C0(n500), 
        .C1(addrD[1]), .Y(n497) );
  AOI31 U565 ( .A0(n501), .A1(n502), .A2(n503), .B0(n504), .Y(n496) );
  NOR2B U566 ( .AN(n505), .B(n506), .Y(n503) );
  NOR4B U567 ( .AN(n507), .B(n508), .C(n509), .D(n510), .Y(n494) );
  OAI2BB2 U568 ( .B0(n511), .B1(n512), .A0N(n513), .A1N(n514), .Y(n510) );
  OAI32 U569 ( .A0(n515), .A1(n516), .A2(n517), .B0(n518), .B1(n519), .Y(n509)
         );
  NOR2B U570 ( .AN(n520), .B(n521), .Y(n518) );
  AOI31 U571 ( .A0(n522), .A1(n523), .A2(n524), .B0(n525), .Y(n507) );
  NAND2B U572 ( .AN(n526), .B(n527), .Y(n701) );
  AOI222 U573 ( .A0(db_o[0]), .A1(n458), .B0(n500), .B1(addrD[0]), .C0(n528), 
        .C1(n529), .Y(n527) );
  OAI222 U574 ( .A0(n530), .A1(n495), .B0(n531), .B1(n532), .C0(n533), .C1(
        n487), .Y(n526) );
  AOI21 U575 ( .A0(n511), .A1(n534), .B0(n514), .Y(n531) );
  NOR3B U576 ( .AN(addrT[4]), .B(n535), .C(n520), .Y(n514) );
  AOI211 U577 ( .A0(n536), .A1(n537), .B0(n538), .C0(n508), .Y(n530) );
  OAI221 U578 ( .A0(n502), .A1(n539), .B0(addrT[3]), .B1(n540), .C0(n541), .Y(
        n508) );
  OR2 U579 ( .A(n520), .B(n542), .Y(n539) );
  OAI33 U580 ( .A0(n519), .A1(n543), .A2(n520), .B0(n544), .B1(addrT[3]), .B2(
        n545), .Y(n538) );
  NOR2B U581 ( .AN(n505), .B(addrT[0]), .Y(n543) );
  INV U582 ( .A(n546), .Y(n702) );
  AOI221 U583 ( .A0(db_o[7]), .A1(n458), .B0(n547), .B1(n548), .C0(n499), .Y(
        n546) );
  OAI211 U584 ( .A0(n549), .A1(n550), .B0(n551), .C0(n552), .Y(n548) );
  AOI221 U585 ( .A0(addrT[3]), .A1(n553), .B0(n554), .B1(n555), .C0(n556), .Y(
        n552) );
  NOR2B U586 ( .AN(n521), .B(addrT[1]), .Y(n554) );
  OAI21 U587 ( .A0(n545), .A1(n557), .B0(n558), .Y(n553) );
  INV U588 ( .A(\decider/N64 ), .Y(n703) );
  INV U589 ( .A(\decider/N63 ), .Y(n704) );
  INV U590 ( .A(\decider/N62 ), .Y(n705) );
  INV U591 ( .A(\decider/N61 ), .Y(n706) );
  INV U592 ( .A(\decider/N60 ), .Y(n707) );
  INV U593 ( .A(\r62/PROD1[4] ), .Y(n708) );
  INV U594 ( .A(\decider/N58 ), .Y(n709) );
  INV U595 ( .A(\decider/N57 ), .Y(n710) );
  OAI21 U596 ( .A0(\decider/posy_m_rex_top[9] ), .A1(n451), .B0(n560), .Y(n713) );
  OAI21 U597 ( .A0(\decider/posy_m_rex_top[8] ), .A1(n451), .B0(n560), .Y(n714) );
  OAI21 U598 ( .A0(\decider/posy_m_rex_top[7] ), .A1(n451), .B0(n560), .Y(n715) );
  OAI21 U599 ( .A0(\decider/posy_m_rex_top[6] ), .A1(n451), .B0(n560), .Y(n716) );
  INV U600 ( .A(n561), .Y(n717) );
  MX2 U601 ( .A(\decider/posy_m_obstacle_top [5]), .B(
        \decider/posy_m_rex_top[5] ), .S0(n452), .Y(n561) );
  INV U602 ( .A(n562), .Y(n718) );
  MX2 U603 ( .A(\decider/posy_m_obstacle_top [4]), .B(
        \decider/posy_m_rex_top[4] ), .S0(n453), .Y(n562) );
  INV U604 ( .A(n563), .Y(n719) );
  MX2 U605 ( .A(\decider/posy_m_obstacle_top [3]), .B(
        \decider/posy_m_rex_top[3] ), .S0(n454), .Y(n563) );
  INV U606 ( .A(n564), .Y(n720) );
  MX2 U607 ( .A(addrD[2]), .B(\decider/posy_m_rex_top[2] ), .S0(n455), .Y(n564) );
  OAI21 U608 ( .A0(\decider/posy_m_rex_top[14] ), .A1(n451), .B0(n560), .Y(
        n722) );
  OAI21 U609 ( .A0(\decider/posy_m_rex_top[13] ), .A1(n451), .B0(n560), .Y(
        n723) );
  OAI21 U610 ( .A0(\decider/posy_m_rex_top[12] ), .A1(n451), .B0(n560), .Y(
        n724) );
  OAI21 U611 ( .A0(\decider/posy_m_rex_top[11] ), .A1(n451), .B0(n560), .Y(
        n725) );
  OAI21 U612 ( .A0(\decider/posy_m_rex_top[10] ), .A1(n451), .B0(n560), .Y(
        n726) );
  INV U613 ( .A(n721), .Y(n560) );
  NOR2B U614 ( .AN(n406), .B(n451), .Y(n721) );
  INV U615 ( .A(n565), .Y(n727) );
  MX2 U616 ( .A(n732), .B(\decider/posy_m_rex_top[1] ), .S0(n452), .Y(n565) );
  MX2 U617 ( .A(addrD[0]), .B(\decider/rex_top [0]), .S0(n453), .Y(n728) );
  INV U618 ( .A(addrD[1]), .Y(n732) );
  MX2 U619 ( .A(n566), .B(n567), .S0(addrD[5]), .Y(n398) );
  OAI21 U620 ( .A0(addrD[4]), .A1(n568), .B0(n569), .Y(n567) );
  NOR2B U621 ( .AN(n570), .B(n568), .Y(n566) );
  MX2 U622 ( .A(n571), .B(n572), .S0(addrD[0]), .Y(n397) );
  MX2 U623 ( .A(n573), .B(n574), .S0(addrD[1]), .Y(n396) );
  INV U624 ( .A(n575), .Y(n574) );
  NOR2B U625 ( .AN(addrD[0]), .B(n568), .Y(n573) );
  MX2 U626 ( .A(n576), .B(n577), .S0(addrD[2]), .Y(n395) );
  OAI21 U627 ( .A0(addrD[1]), .A1(n568), .B0(n575), .Y(n577) );
  AOI2BB1 U628 ( .A0N(addrD[0]), .A1N(n568), .B0(n572), .Y(n575) );
  NOR3B U629 ( .AN(addrD[1]), .B(n568), .C(n731), .Y(n576) );
  MX2 U630 ( .A(n578), .B(n579), .S0(addrD[3]), .Y(n394) );
  NOR2B U631 ( .AN(n580), .B(n568), .Y(n578) );
  MX2 U632 ( .A(n581), .B(n582), .S0(addrD[4]), .Y(n393) );
  INV U633 ( .A(n569), .Y(n582) );
  AOI2BB1 U634 ( .A0N(addrD[3]), .A1N(n568), .B0(n579), .Y(n569) );
  OAI21 U635 ( .A0(n580), .A1(n568), .B0(n583), .Y(n579) );
  NOR3B U636 ( .AN(n580), .B(n568), .C(n734), .Y(n581) );
  OAI2BB2 U637 ( .B0(n584), .B1(n585), .A0N(\driver/N47 ), .A1N(n446), .Y(n392) );
  MX2 U638 ( .A(n446), .B(n587), .S0(addrD[6]), .Y(n391) );
  OAI2BB2 U639 ( .B0(n588), .B1(n584), .A0N(\driver/N44 ), .A1N(n446), .Y(n390) );
  OAI2BB2 U640 ( .B0(n584), .B1(n589), .A0N(\driver/N45 ), .A1N(n446), .Y(n389) );
  OAI2BB2 U641 ( .B0(n584), .B1(n590), .A0N(\driver/N46 ), .A1N(n446), .Y(n388) );
  NOR3B U642 ( .AN(n448), .B(n587), .C(\driver/N17 ), .Y(n586) );
  OAI21 U643 ( .A0(n729), .A1(n591), .B0(n592), .Y(n387) );
  NAND2 U644 ( .A(n593), .B(n592), .Y(n386) );
  MX2 U645 ( .A(n594), .B(n595), .S0(n596), .Y(n593) );
  AOI31 U646 ( .A0(cs_o[3]), .A1(addrD[8]), .A2(n597), .B0(n598), .Y(n594) );
  NOR3B U647 ( .AN(n448), .B(n487), .C(n588), .Y(n597) );
  INV U648 ( .A(addrD[7]), .Y(n588) );
  OAI31 U649 ( .A0(n599), .A1(n600), .A2(n583), .B0(n568), .Y(n385) );
  INV U650 ( .A(n571), .Y(n568) );
  NOR3B U651 ( .AN(n448), .B(n572), .C(\driver/N17 ), .Y(n571) );
  INV U652 ( .A(n572), .Y(n583) );
  AOI21 U653 ( .A0(en_o), .A1(n601), .B0(n602), .Y(n572) );
  INV U654 ( .A(dori_o), .Y(n599) );
  INV U655 ( .A(n603), .Y(n384) );
  AOI222 U656 ( .A0(n457), .A1(\decider/N87 ), .B0(addrT[0]), .B1(n449), .C0(
        n453), .C1(\decider/N86 ), .Y(n603) );
  INV U657 ( .A(n605), .Y(n383) );
  AOI222 U658 ( .A0(n457), .A1(\decider/N88 ), .B0(addrT[1]), .B1(n449), .C0(
        n452), .C1(\decider/N85 ), .Y(n605) );
  INV U659 ( .A(n606), .Y(n382) );
  AOI222 U660 ( .A0(n457), .A1(\decider/N89 ), .B0(addrT[2]), .B1(n449), .C0(
        n455), .C1(\decider/N84 ), .Y(n606) );
  INV U661 ( .A(n607), .Y(n381) );
  AOI222 U662 ( .A0(n457), .A1(\decider/N90 ), .B0(addrT[3]), .B1(n449), .C0(
        n454), .C1(\decider/N83 ), .Y(n607) );
  INV U663 ( .A(n608), .Y(n380) );
  AOI222 U664 ( .A0(n457), .A1(\decider/N91 ), .B0(addrT[4]), .B1(n449), .C0(
        n453), .C1(\decider/N82 ), .Y(n608) );
  INV U665 ( .A(n609), .Y(n379) );
  AOI222 U666 ( .A0(n457), .A1(\decider/N92 ), .B0(addrT[5]), .B1(n449), .C0(
        n452), .C1(\decider/N81 ), .Y(n609) );
  INV U667 ( .A(n610), .Y(n378) );
  AOI222 U668 ( .A0(n457), .A1(\decider/N93 ), .B0(addrT[6]), .B1(n449), .C0(
        n455), .C1(\decider/N80 ), .Y(n610) );
  INV U669 ( .A(n611), .Y(n377) );
  AOI222 U670 ( .A0(n457), .A1(\decider/N94 ), .B0(addrT[7]), .B1(n449), .C0(
        n454), .C1(\decider/N79 ), .Y(n611) );
  INV U671 ( .A(n612), .Y(n376) );
  AOI222 U672 ( .A0(n457), .A1(\decider/N95 ), .B0(n449), .B1(addrT[8]), .C0(
        n453), .C1(\decider/N78 ), .Y(n612) );
  INV U673 ( .A(n613), .Y(n375) );
  AOI222 U674 ( .A0(n457), .A1(\decider/N96 ), .B0(n449), .B1(addrT[9]), .C0(
        n452), .C1(\decider/N77 ), .Y(n613) );
  NOR3B U675 ( .AN(n451), .B(n435), .C(\decider/obstacle_right [15]), .Y(n604)
         );
  NOR2B U676 ( .AN(n406), .B(\decider/sub_75/carry[6] ), .Y(n559) );
  INV U677 ( .A(n614), .Y(n372) );
  AOI221 U678 ( .A0(n500), .A1(addrD[2]), .B0(db_o[2]), .B1(n458), .C0(n615), 
        .Y(n614) );
  OAI221 U679 ( .A0(n616), .A1(n495), .B0(n533), .B1(n589), .C0(n617), .Y(n615) );
  INV U680 ( .A(addrD[8]), .Y(n589) );
  AOI211 U681 ( .A0(n556), .A1(n618), .B0(n619), .C0(n620), .Y(n616) );
  OAI211 U682 ( .A0(n621), .A1(n523), .B0(n512), .C0(n622), .Y(n619) );
  INV U683 ( .A(n623), .Y(n622) );
  INV U684 ( .A(n536), .Y(n512) );
  NOR2B U685 ( .AN(n624), .B(addrT[2]), .Y(n536) );
  AOI32 U686 ( .A0(n505), .A1(n502), .A2(n522), .B0(n625), .B1(addrT[1]), .Y(
        n621) );
  NOR2B U687 ( .AN(n626), .B(n515), .Y(n556) );
  INV U688 ( .A(n627), .Y(n371) );
  AOI211 U689 ( .A0(db_o[3]), .A1(n458), .B0(n628), .C0(n629), .Y(n627) );
  OAI222 U690 ( .A0(n630), .A1(n495), .B0(n631), .B1(n532), .C0(n734), .C1(
        n632), .Y(n628) );
  AOI2BB2 U691 ( .B0(n625), .B1(n511), .A0N(n544), .A1N(n524), .Y(n631) );
  INV U692 ( .A(n545), .Y(n524) );
  NOR2B U693 ( .AN(n511), .B(n618), .Y(n545) );
  INV U694 ( .A(n633), .Y(n544) );
  NOR4BB U695 ( .AN(n634), .BN(n635), .C(n624), .D(n636), .Y(n630) );
  AOI31 U696 ( .A0(n535), .A1(n618), .A2(n637), .B0(n638), .Y(n635) );
  AOI221 U697 ( .A0(n639), .A1(n537), .B0(n513), .B1(n623), .C0(n620), .Y(n634) );
  OAI221 U698 ( .A0(n640), .A1(n541), .B0(addrT[3]), .B1(n641), .C0(n642), .Y(
        n620) );
  NOR2 U699 ( .A(n643), .B(n525), .Y(n642) );
  INV U700 ( .A(n637), .Y(n641) );
  OR3 U701 ( .A(n520), .B(n523), .C(n618), .Y(n541) );
  AOI2BB2 U702 ( .B0(addrT[4]), .B1(n549), .A0N(n537), .A1N(addrT[6]), .Y(n640) );
  INV U703 ( .A(n644), .Y(n370) );
  AOI211 U704 ( .A0(db_o[4]), .A1(n458), .B0(n645), .C0(n629), .Y(n644) );
  OAI222 U705 ( .A0(n646), .A1(n495), .B0(n647), .B1(n532), .C0(n735), .C1(
        n632), .Y(n645) );
  AOI2BB2 U706 ( .B0(n648), .B1(addrT[2]), .A0N(addrT[1]), .A1N(n540), .Y(n647) );
  NOR4 U707 ( .A(n636), .B(n649), .C(n525), .D(n643), .Y(n646) );
  OAI21 U708 ( .A0(n517), .A1(n650), .B0(n651), .Y(n649) );
  AOI33 U709 ( .A0(n624), .A1(n523), .A2(addrT[1]), .B0(n521), .B1(n652), .B2(
        n653), .Y(n651) );
  OAI31 U710 ( .A0(n618), .A1(n511), .A2(n502), .B0(n654), .Y(n653) );
  AOI211 U711 ( .A0(n513), .A1(n655), .B0(n656), .C0(n624), .Y(n650) );
  OAI221 U712 ( .A0(n657), .A1(n495), .B0(n730), .B1(n632), .C0(n658), .Y(n369) );
  AOI21 U713 ( .A0(db_o[5]), .A1(n458), .B0(n629), .Y(n658) );
  NAND2B U714 ( .AN(n504), .B(n533), .Y(n629) );
  INV U715 ( .A(n499), .Y(n533) );
  NOR2B U716 ( .AN(n659), .B(n660), .Y(n499) );
  INV U717 ( .A(n617), .Y(n504) );
  OAI21 U718 ( .A0(n601), .A1(n528), .B0(n529), .Y(n617) );
  INV U719 ( .A(addrD[5]), .Y(n730) );
  NOR3B U720 ( .AN(n661), .B(n662), .C(n663), .Y(n657) );
  MX2 U721 ( .A(n636), .B(n664), .S0(addrT[0]), .Y(n663) );
  NOR3B U722 ( .AN(addrT[2]), .B(n550), .C(addrT[1]), .Y(n664) );
  INV U723 ( .A(n626), .Y(n550) );
  NOR2B U724 ( .AN(n623), .B(addrT[1]), .Y(n636) );
  NOR3B U725 ( .AN(n625), .B(addrT[3]), .C(addrT[2]), .Y(n623) );
  NOR2B U726 ( .AN(n534), .B(n502), .Y(n625) );
  AOI221 U727 ( .A0(n665), .A1(n624), .B0(addrT[3]), .B1(n666), .C0(n638), .Y(
        n661) );
  NOR3B U728 ( .AN(n513), .B(n516), .C(n517), .Y(n638) );
  INV U729 ( .A(n665), .Y(n517) );
  OAI221 U730 ( .A0(n549), .A1(n667), .B0(n540), .B1(n515), .C0(n668), .Y(n666) );
  AOI221 U731 ( .A0(n522), .A1(n669), .B0(n670), .B1(n626), .C0(n656), .Y(n668) );
  NOR3B U732 ( .AN(n521), .B(addrT[1]), .C(n502), .Y(n656) );
  NOR2B U733 ( .AN(n671), .B(n502), .Y(n626) );
  NOR2B U734 ( .AN(addrT[1]), .B(addrT[0]), .Y(n670) );
  NAND2B U735 ( .AN(n515), .B(n618), .Y(n669) );
  INV U736 ( .A(n537), .Y(n515) );
  INV U737 ( .A(n624), .Y(n540) );
  INV U738 ( .A(n648), .Y(n667) );
  NOR2B U739 ( .AN(n655), .B(addrT[4]), .Y(n624) );
  OAI211 U740 ( .A0(n672), .A1(n495), .B0(n632), .C0(n673), .Y(n368) );
  AOI2BB2 U741 ( .B0(db_o[6]), .B1(n458), .A0N(n674), .A1N(n532), .Y(n673) );
  INV U742 ( .A(n501), .Y(n532) );
  NOR2B U743 ( .AN(n547), .B(n523), .Y(n501) );
  AOI211 U744 ( .A0(n633), .A1(n675), .B0(n676), .C0(n677), .Y(n674) );
  MX2 U745 ( .A(n648), .B(n678), .S0(n537), .Y(n677) );
  NOR2B U746 ( .AN(n535), .B(addrT[0]), .Y(n537) );
  NOR2B U747 ( .AN(addrT[4]), .B(n506), .Y(n678) );
  OAI31 U748 ( .A0(n513), .A1(addrT[1]), .A2(n557), .B0(n558), .Y(n676) );
  INV U749 ( .A(n522), .Y(n558) );
  INV U750 ( .A(n671), .Y(n557) );
  INV U751 ( .A(n505), .Y(n675) );
  NOR2B U752 ( .AN(addrT[2]), .B(n535), .Y(n505) );
  NOR2B U753 ( .AN(n671), .B(addrT[4]), .Y(n633) );
  INV U754 ( .A(n500), .Y(n632) );
  NOR2B U755 ( .AN(n598), .B(n660), .Y(n500) );
  INV U756 ( .A(n529), .Y(n660) );
  INV U757 ( .A(n547), .Y(n495) );
  NOR4 U758 ( .A(addrT[9]), .B(addrT[8]), .C(\r62/ab[12][2] ), .D(n679), .Y(
        n547) );
  OAI211 U759 ( .A0(n680), .A1(n455), .B0(n448), .C0(n529), .Y(n679) );
  NOR2B U760 ( .AN(rstn), .B(n458), .Y(n529) );
  AOI211 U761 ( .A0(en_o), .A1(n681), .B0(n600), .C0(n602), .Y(n498) );
  OAI2BB1 U762 ( .A0N(en_o), .A1N(n448), .B0(rstn), .Y(n602) );
  NOR2 U763 ( .A(n435), .B(\decider/sub_75/carry[6] ), .Y(n680) );
  AOI31 U764 ( .A0(n671), .A1(n513), .A2(n665), .B0(n662), .Y(n672) );
  OAI211 U765 ( .A0(n654), .A1(n506), .B0(n551), .C0(n682), .Y(n662) );
  AOI21 U766 ( .A0(addrT[2]), .A1(n683), .B0(n643), .Y(n682) );
  NOR2B U767 ( .AN(n639), .B(n549), .Y(n643) );
  OAI2BB2 U768 ( .B0(n506), .B1(n519), .A0N(addrT[3]), .A1N(n648), .Y(n683) );
  NOR2B U769 ( .AN(n534), .B(addrT[4]), .Y(n648) );
  NOR2B U770 ( .AN(n542), .B(n520), .Y(n534) );
  NAND2B U771 ( .AN(addrT[7]), .B(n652), .Y(n520) );
  INV U772 ( .A(addrT[6]), .Y(n542) );
  NOR3 U773 ( .A(n637), .B(n525), .C(n684), .Y(n551) );
  NOR4BB U774 ( .AN(addrT[7]), .BN(n555), .C(addrT[6]), .D(n511), .Y(n684) );
  NOR4BB U775 ( .AN(n523), .BN(n618), .C(addrT[5]), .D(addrT[4]), .Y(n555) );
  NOR2B U776 ( .AN(n639), .B(n618), .Y(n525) );
  NOR2B U777 ( .AN(n523), .B(n516), .Y(n639) );
  INV U778 ( .A(n655), .Y(n516) );
  NOR2B U779 ( .AN(n671), .B(addrT[6]), .Y(n655) );
  NOR2B U780 ( .AN(n522), .B(n502), .Y(n637) );
  INV U781 ( .A(addrT[4]), .Y(n502) );
  NOR2B U782 ( .AN(n521), .B(n652), .Y(n522) );
  INV U783 ( .A(addrT[5]), .Y(n652) );
  INV U784 ( .A(n521), .Y(n506) );
  NOR2B U785 ( .AN(addrT[6]), .B(addrT[7]), .Y(n521) );
  AOI2BB2 U786 ( .B0(addrT[4]), .B1(n665), .A0N(n549), .A1N(n519), .Y(n654) );
  NAND2B U787 ( .AN(addrT[3]), .B(addrT[4]), .Y(n519) );
  INV U788 ( .A(n511), .Y(n549) );
  NOR2B U789 ( .AN(addrT[0]), .B(n535), .Y(n511) );
  INV U790 ( .A(addrT[1]), .Y(n535) );
  NOR2B U791 ( .AN(n618), .B(n523), .Y(n665) );
  INV U792 ( .A(addrT[3]), .Y(n523) );
  INV U793 ( .A(addrT[2]), .Y(n618) );
  INV U794 ( .A(addrT[0]), .Y(n513) );
  NOR2B U795 ( .AN(addrT[5]), .B(addrT[7]), .Y(n671) );
  NOR2B U796 ( .AN(n592), .B(n681), .Y(n367) );
  OAI31 U797 ( .A0(n685), .A1(\driver/N17 ), .A2(n528), .B0(n729), .Y(n592) );
  INV U798 ( .A(n596), .Y(n729) );
  AOI211 U799 ( .A0(en_o), .A1(n685), .B0(n600), .C0(n584), .Y(n596) );
  INV U800 ( .A(n587), .Y(n584) );
  AOI2BB1 U801 ( .A0N(n686), .A1N(n687), .B0(\driver/N17 ), .Y(n587) );
  AOI31 U802 ( .A0(n570), .A1(addrD[5]), .A2(n448), .B0(n601), .Y(n687) );
  NOR3B U803 ( .AN(n681), .B(n688), .C(start), .Y(n601) );
  INV U804 ( .A(\driver/start_history [1]), .Y(n688) );
  NOR2B U805 ( .AN(n689), .B(n591), .Y(n681) );
  INV U806 ( .A(state[2]), .Y(n591) );
  NOR3B U807 ( .AN(n580), .B(n734), .C(n735), .Y(n570) );
  INV U808 ( .A(addrD[4]), .Y(n735) );
  INV U809 ( .A(addrD[3]), .Y(n734) );
  NOR3B U810 ( .AN(addrD[1]), .B(n731), .C(n733), .Y(n580) );
  INV U811 ( .A(addrD[2]), .Y(n733) );
  INV U812 ( .A(addrD[0]), .Y(n731) );
  INV U813 ( .A(en_o), .Y(n686) );
  INV U814 ( .A(n690), .Y(n600) );
  OAI31 U815 ( .A0(n659), .A1(n528), .A2(n598), .B0(en_o), .Y(n690) );
  NOR3B U816 ( .AN(state[1]), .B(state[0]), .C(state[2]), .Y(n598) );
  NOR3B U817 ( .AN(state[0]), .B(state[2]), .C(state[1]), .Y(n659) );
  NOR2B U818 ( .AN(n689), .B(state[2]), .Y(n528) );
  NOR2B U819 ( .AN(state[2]), .B(n689), .Y(n685) );
  NOR2B U820 ( .AN(state[1]), .B(n595), .Y(n689) );
  NOR3B U821 ( .AN(n595), .B(state[2]), .C(state[1]), .Y(n366) );
  INV U822 ( .A(state[0]), .Y(n595) );
  XOR2 U823 ( .A(n691), .B(start), .Y(n356) );
  NOR2B U824 ( .AN(rstn), .B(en_o), .Y(\driver/N96 ) );
  INV U825 ( .A(rstn), .Y(\driver/N17 ) );
  NOR2B U826 ( .AN(addrD[10]), .B(n590), .Y(cs_o[3]) );
  NOR2B U827 ( .AN(addrD[10]), .B(addrD[9]), .Y(cs_o[2]) );
  NOR2B U828 ( .AN(n585), .B(n590), .Y(cs_o[1]) );
  INV U829 ( .A(addrD[9]), .Y(n590) );
  NOR2B U830 ( .AN(\clock_divider/N17 ), .B(n691), .Y(\clock_divider/N30 ) );
  NOR2B U831 ( .AN(\clock_divider/N16 ), .B(n691), .Y(\clock_divider/N29 ) );
  NOR2B U832 ( .AN(\clock_divider/N15 ), .B(n691), .Y(\clock_divider/N28 ) );
  NOR2B U833 ( .AN(\clock_divider/N14 ), .B(n691), .Y(\clock_divider/N27 ) );
  NOR2B U834 ( .AN(\clock_divider/N13 ), .B(n691), .Y(\clock_divider/N26 ) );
  NOR2B U835 ( .AN(\clock_divider/N12 ), .B(n691), .Y(\clock_divider/N25 ) );
  NOR2B U836 ( .AN(\clock_divider/N11 ), .B(n691), .Y(\clock_divider/N24 ) );
  NOR2B U837 ( .AN(\clock_divider/N10 ), .B(n691), .Y(\clock_divider/N23 ) );
  NOR2B U838 ( .AN(\clock_divider/N9 ), .B(n691), .Y(\clock_divider/N22 ) );
  NOR2B U839 ( .AN(\clock_divider/N8 ), .B(n691), .Y(\clock_divider/N21 ) );
  NOR2B U840 ( .AN(\clock_divider/N7 ), .B(n691), .Y(\clock_divider/N20 ) );
  NOR2B U841 ( .AN(\clock_divider/N6 ), .B(n691), .Y(\clock_divider/N19 ) );
  AND2 U842 ( .A(n692), .B(n693), .Y(n691) );
  NOR4BB U843 ( .AN(n694), .BN(\clock_divider/cnt5k[0] ), .C(
        \clock_divider/cnt5k[11] ), .D(\clock_divider/cnt5k[10] ), .Y(n693) );
  NOR4 U844 ( .A(\clock_divider/cnt5k[6] ), .B(\clock_divider/cnt5k[5] ), .C(
        \clock_divider/cnt5k[4] ), .D(\clock_divider/cnt5k[3] ), .Y(n694) );
  AND4 U845 ( .A(\clock_divider/cnt5k[8] ), .B(\clock_divider/cnt5k[7] ), .C(
        \clock_divider/cnt5k[9] ), .D(n695), .Y(n692) );
  AND3 U846 ( .A(\clock_divider/cnt5k[1] ), .B(\clock_divider/cnt5k[12] ), .C(
        \clock_divider/cnt5k[2] ), .Y(n695) );
  INV U847 ( .A(\clock_divider/cnt5k[0] ), .Y(\clock_divider/N18 ) );
  MX2 U848 ( .A(\decider/N77 ), .B(\decider/N64 ), .S0(n454), .Y(\U1/U5/Z_9 )
         );
  MX2 U849 ( .A(\decider/N78 ), .B(\decider/N63 ), .S0(n455), .Y(\U1/U5/Z_8 )
         );
  MX2 U850 ( .A(\decider/N79 ), .B(\decider/N62 ), .S0(n452), .Y(\U1/U5/Z_7 )
         );
  MX2 U851 ( .A(\decider/N80 ), .B(\decider/N61 ), .S0(n453), .Y(\U1/U5/Z_6 )
         );
  MX2 U852 ( .A(\decider/N81 ), .B(\decider/N60 ), .S0(n454), .Y(\U1/U5/Z_5 )
         );
  MX2 U853 ( .A(\decider/N82 ), .B(\r62/PROD1[4] ), .S0(n455), .Y(\U1/U5/Z_4 )
         );
  MX2 U854 ( .A(\decider/N83 ), .B(\decider/N58 ), .S0(n452), .Y(\U1/U5/Z_3 )
         );
  MX2 U855 ( .A(\decider/N84 ), .B(\decider/N57 ), .S0(n453), .Y(\U1/U5/Z_2 )
         );
  MX2 U856 ( .A(\decider/N71 ), .B(n696), .S0(n454), .Y(\U1/U5/Z_15 ) );
  MX2 U857 ( .A(\decider/N72 ), .B(n697), .S0(n455), .Y(\U1/U5/Z_14 ) );
  MX2 U858 ( .A(\decider/N73 ), .B(\r62/A1[11] ), .S0(n452), .Y(\U1/U5/Z_13 )
         );
  MX2 U859 ( .A(\decider/N74 ), .B(\r62/SUMB[12][0] ), .S0(n453), .Y(
        \U1/U5/Z_12 ) );
  MX2 U860 ( .A(\decider/N75 ), .B(\r62/A1[9] ), .S0(n454), .Y(\U1/U5/Z_11 )
         );
  MX2 U861 ( .A(\decider/N76 ), .B(\decider/N65 ), .S0(n455), .Y(\U1/U5/Z_10 )
         );
  OAI2BB1 U862 ( .A0N(n406), .A1N(\decider/N85 ), .B0(n711), .Y(\U1/U5/Z_1 )
         );
  NAND2B U863 ( .AN(n406), .B(\U1/U3/Z_1 ), .Y(n711) );
  OAI2BB1 U864 ( .A0N(n406), .A1N(\decider/N86 ), .B0(n712), .Y(\U1/U5/Z_0 )
         );
  NAND2B U865 ( .AN(n406), .B(\U1/U3/Z_0 ), .Y(n712) );
  NOR2B U866 ( .AN(\decider/obstacle_right [12]), .B(n452), .Y(\r62/ab[9][2] )
         );
  NOR2B U867 ( .AN(\decider/obstacle_right [11]), .B(n453), .Y(\r62/ab[8][2] )
         );
  NOR2B U868 ( .AN(\decider/obstacle_right [10]), .B(n454), .Y(\r62/ab[7][2] )
         );
  NOR2B U869 ( .AN(\decider/obstacle_right [9]), .B(n455), .Y(\r62/ab[6][2] )
         );
  NOR2B U870 ( .AN(\decider/obstacle_right [8]), .B(n452), .Y(\r62/ab[5][2] )
         );
  MX2 U871 ( .A(\decider/obstacle_right [7]), .B(\decider/posx_m_rex_left [7]), 
        .S0(n452), .Y(\U1/U3/Z_4 ) );
  MX2 U872 ( .A(\decider/obstacle_right [6]), .B(\decider/posx_m_rex_left [6]), 
        .S0(n453), .Y(\U1/U3/Z_3 ) );
  MX2 U873 ( .A(\decider/obstacle_right [5]), .B(\decider/posx_m_rex_left [5]), 
        .S0(n454), .Y(\U1/U3/Z_2 ) );
  NOR2B U874 ( .AN(\decider/obstacle_right [15]), .B(n453), .Y(\r62/ab[12][2] ) );
  NOR2B U875 ( .AN(\decider/obstacle_right [14]), .B(n454), .Y(\r62/ab[11][2] ) );
  NOR2B U876 ( .AN(\decider/obstacle_right [13]), .B(n455), .Y(\r62/ab[10][2] ) );
  MX2 U877 ( .A(\decider/obstacle_right [4]), .B(\decider/posx_m_rex_left [4]), 
        .S0(n455), .Y(\U1/U3/Z_1 ) );
  MX2 U878 ( .A(\decider/obstacle_right [3]), .B(n487), .S0(n452), .Y(
        \U1/U3/Z_0 ) );
  MX2 U879 ( .A(n696), .B(\decider/N102 ), .S0(n453), .Y(\U1/U2/Z_15 ) );
  XOR2 U880 ( .A(\r62/A1[13] ), .B(n698), .Y(n696) );
  AND2 U881 ( .A(n428), .B(\r62/SUMB[12][2] ), .Y(n698) );
  MX2 U882 ( .A(n697), .B(\decider/N101 ), .S0(n454), .Y(\U1/U2/Z_14 ) );
  XOR2 U883 ( .A(\r62/SUMB[12][2] ), .B(n428), .Y(n697) );
  MX2 U884 ( .A(\r62/A1[11] ), .B(\decider/N100 ), .S0(n455), .Y(\U1/U2/Z_13 )
         );
  MX2 U885 ( .A(\r62/SUMB[12][0] ), .B(\decider/N99 ), .S0(n452), .Y(
        \U1/U2/Z_12 ) );
  MX2 U886 ( .A(\r62/A1[9] ), .B(\decider/N98 ), .S0(n453), .Y(\U1/U2/Z_11 )
         );
  MX2 U887 ( .A(\decider/N65 ), .B(\decider/N97 ), .S0(n454), .Y(\U1/U2/Z_10 )
         );
  NOR2 U888 ( .A(addrD[8]), .B(\decider/rex_top [15]), .Y(n699) );
  NOR2B U889 ( .AN(n585), .B(addrD[9]), .Y(cs_o[0]) );
  INV U890 ( .A(addrD[10]), .Y(n585) );
  GameCenter gamecenter ( .clk(clk), .rstn(rstn), .in_up(jmp_key), .rex_y(
        rex_down), .obstacle_x(obstacle_left) );
endmodule

