
module FDE_Rex_Runner ( clk, rstn, db_o, dori_o, cs_o, en_o, rw_o, rst_o, 
        state );
  output [7:0] db_o;
  output [3:0] cs_o;
  output [2:0] state;
  input clk, rstn;
  output dori_o, en_o, rw_o, rst_o;
  wire   start, \driver/N96 , \driver/N47 , \driver/N46 , \driver/N45 ,
         \driver/N44 , \driver/*Logic0* , \decider/N96 , \decider/N95 ,
         \decider/N94 , \decider/N93 , \decider/N92 , \decider/N91 ,
         \decider/N90 , \decider/N89 , \decider/N88 , \decider/N85 ,
         \decider/N84 , \decider/N83 , \decider/N82 , \decider/N81 ,
         \decider/N80 , \decider/N79 , \decider/N78 , \decider/N77 ,
         \decider/N64 , \decider/N63 , \decider/N62 , \decider/N61 ,
         \decider/N60 , \decider/N58 , \decider/N57 , \decider/N55 ,
         \decider/N38 , \decider/posx_m_obstacle_right[15] ,
         \decider/posy_m_rex_top[1] , \decider/posy_m_rex_top[2] ,
         \decider/posy_m_rex_top[3] , \decider/posy_m_rex_top[4] ,
         \decider/posy_m_rex_top[5] , \clock_divider/N30 , \clock_divider/N29 ,
         \clock_divider/N28 , \clock_divider/N27 , \clock_divider/N26 ,
         \clock_divider/N25 , \clock_divider/N24 , \clock_divider/N23 ,
         \clock_divider/N22 , \clock_divider/N21 , \clock_divider/N20 ,
         \clock_divider/N19 , \clock_divider/N18 , \clock_divider/N17 ,
         \clock_divider/N16 , \clock_divider/N15 , \clock_divider/N14 ,
         \clock_divider/N13 , \clock_divider/N12 , \clock_divider/N11 ,
         \clock_divider/N10 , \clock_divider/N9 , \clock_divider/N8 ,
         \clock_divider/N7 , \clock_divider/N6 , \clock_divider/cnt5k[0] ,
         \clock_divider/cnt5k[1] , \clock_divider/cnt5k[2] ,
         \clock_divider/cnt5k[3] , \clock_divider/cnt5k[4] ,
         \clock_divider/cnt5k[5] , \clock_divider/cnt5k[6] ,
         \clock_divider/cnt5k[7] , \clock_divider/cnt5k[8] ,
         \clock_divider/cnt5k[9] , \clock_divider/cnt5k[10] ,
         \clock_divider/cnt5k[11] , \clock_divider/cnt5k[12] , n329, n330,
         n331, n332, n333, n334, n356, n357, n377, n378, n379, n380, n384,
         n385, n386, n387, n388, n389, n390, n391, n392, n393, n394, n395,
         n396, n397, \r51/carry[9] , \r51/carry[8] , \r51/carry[7] ,
         \r51/carry[6] , \r51/carry[5] , \r51/carry[4] , \r51/carry[3] ,
         \r51/carry[2] , \r51/carry[1] ,
         \add_2_root_decider/add_109_3_cf/carry[2] ,
         \add_2_root_decider/add_109_3_cf/carry[3] ,
         \add_2_root_decider/add_109_3_cf/carry[4] ,
         \add_2_root_decider/add_109_3_cf/carry[6] ,
         \add_2_root_decider/add_109_3_cf/carry[7] , \r62/PROD1[4] ,
         \r62/SUMB[1][2] , \r62/SUMB[1][3] , \r62/SUMB[2][2] ,
         \r62/SUMB[2][3] , \r62/SUMB[3][2] , \r62/SUMB[3][3] ,
         \r62/SUMB[4][2] , \r62/SUMB[4][3] , \r62/SUMB[5][2] ,
         \r62/SUMB[5][3] , \r62/SUMB[6][2] , \r62/SUMB[6][3] ,
         \r62/SUMB[7][2] , \r62/CARRYB[2][2] , \r62/CARRYB[2][3] ,
         \r62/CARRYB[3][0] , \r62/CARRYB[3][2] , \r62/CARRYB[3][3] ,
         \r62/CARRYB[4][0] , \r62/CARRYB[4][2] , \r62/CARRYB[4][3] ,
         \r62/CARRYB[5][2] , \r62/CARRYB[6][2] , \r62/ab[0][2] ,
         \r62/ab[1][0] , \r62/ab[1][2] , \r62/ab[2][0] , \r62/ab[2][2] ,
         \r62/ab[3][0] , \r62/ab[3][2] , \r62/ab[4][0] , \r62/ab[4][2] ,
         \r62/ab[7][2] , \sub_1_root_decider/sub_49/carry[2] ,
         \sub_1_root_decider/sub_49/carry[3] ,
         \sub_1_root_decider/sub_49/carry[5] ,
         \sub_1_root_decider/sub_49/carry[6] , \decider/sub_45/carry[2] ,
         \decider/sub_45/carry[3] , \decider/sub_45/carry[4] ,
         \decider/sub_45/carry[5] , \decider/sub_75/carry[6] ,
         \decider/sub_75/carry[5] , \sub_0_root_decider/sub_73/carry[15] ,
         \r187/carry[8] , \r187/carry[7] , n401, n402, n403, n404, n405, n406,
         n407, n408, n409, n410, n411, n412, n413, n414, n415, n416, n417,
         n418, n419, n420, n421, n422, n423, n424, n425, n426, n427, n428,
         n429, n430, n431, n432, n433, n434, n435, n436, n437, n438, n439,
         n440, n441, n442, n443, n444, n445, n446, n447, n448, n449, n450,
         n451, n452, n453, n454, n455, n456, n457, n458, n459, n460, n461,
         n462, n463, n464, n465, n466, n467, n468, n469, n470, n471, n472,
         n473, n474, n475, n476, n477, n478, n479, n480, n481, n482, n483,
         n484, n485, n486, n487, n488, n489, n490, n491, n492, n493, n494,
         n495, n496, n497, n498, n499, n500, n501, n502, n503, n504, n505,
         n506, n507, n508, n509, n510, n511, n512, n513, n514, n515, n516,
         n517, n518, n519, n520, n521, n522, n523, n524, n525, n526, n527,
         n528, n529, n530, n531, n532, n533, n534, n535, n536, n537, n538,
         n539, n540, n541, n542, n543, n544, n545, n546, n547, n548, n549,
         n550, n551, n552, n553, n554, n555, n556, n557, n558, n559, n560,
         n561, n562, n563, n564, n565, n566, n567, n568, n569, n570, n571,
         n572, n573, n574, n575, n576, n577, n578, n579, n580, n581, n582,
         n583, n584, n585, n586, n587, n588, n589, n590, n591, n592, n593,
         n594, n595, n596, n597, n598, n599, n600, n601, n602, n603, n604,
         n605, n606, n607, n608, n609, n610, n611, n612, n613, n614, n615,
         n616, n617, n618, n619, n620, n621, n622, n623, n624, n625, n626,
         n627, n628, n629, n630, n631, n632, n633, n634, n635, n636, n637,
         n638, n639, n640, n641, n642, n643, n644, n645, n646, n647, n648,
         n649, n650, n651, n652, n653, n654, n655, n656, n657, n658, n659,
         n660, n661, n662, n663, n664, n665, n666, n667, n668, n669, n670,
         n671, n672, n673, n674, n675, n676, n677, n678, n679, n680, n681,
         n682;
  wire   [10:0] addrD;
  wire   [15:0] addrT;
  wire   [1:0] \driver/start_history ;
  wire   [5:0] \decider/posy_m_obstacle_top ;
  wire   [15:0] \decider/obstacle_right ;
  wire   [7:3] \decider/posx_m_rex_left ;
  assign rw_o = \driver/*Logic0* ;

  DFFHQ \driver/en_o_reg  ( .D(\driver/N96 ), .CK(clk), .Q(en_o) );
  DFFHQ \driver/rst_o_reg  ( .D(n649), .CK(clk), .Q(rst_o) );
  DFFRHQ \clock_divider/cnt5k_reg[12]  ( .D(\clock_divider/N30 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[12] ) );
  DFFRHQ \clock_divider/clk_12Hz_reg  ( .D(n356), .CK(clk), .RN(rstn), .Q(
        start) );
  EDFFHQ \driver/start_history_reg[0]  ( .D(start), .E(rstn), .CK(clk), .Q(
        \driver/start_history [0]) );
  EDFFHQ \driver/start_history_reg[1]  ( .D(\driver/start_history [0]), .E(
        rstn), .CK(clk), .Q(\driver/start_history [1]) );
  DFFHQ \driver/y_reg[4]  ( .D(n392), .CK(clk), .Q(addrD[4]) );
  DFFHQ \driver/x_reg[4]  ( .D(n391), .CK(clk), .Q(addrD[10]) );
  DFFHQ \driver/x_reg[0]  ( .D(n390), .CK(clk), .Q(addrD[6]) );
  DFFHQ \driver/x_reg[1]  ( .D(n389), .CK(clk), .Q(addrD[7]) );
  DFFHQ \driver/x_reg[2]  ( .D(n388), .CK(clk), .Q(addrD[8]) );
  DFFHQ \driver/x_reg[3]  ( .D(n387), .CK(clk), .Q(addrD[9]) );
  DFFHQ \driver/state_reg[0]  ( .D(n385), .CK(clk), .Q(state[0]) );
  DFFHQ \driver/state_reg[1]  ( .D(n384), .CK(clk), .Q(state[1]) );
  DFFHQ \driver/state_reg[2]  ( .D(n386), .CK(clk), .Q(state[2]) );
  DFFHQ \driver/y_reg[5]  ( .D(n397), .CK(clk), .Q(addrD[5]) );
  DFFHQ \driver/y_reg[0]  ( .D(n396), .CK(clk), .Q(addrD[0]) );
  DFFHQ \driver/y_reg[1]  ( .D(n395), .CK(clk), .Q(addrD[1]) );
  DFFHQ \driver/y_reg[2]  ( .D(n394), .CK(clk), .Q(addrD[2]) );
  DFFHQ \driver/y_reg[3]  ( .D(n393), .CK(clk), .Q(addrD[3]) );
  DFFHQ \driver/dori_o_reg  ( .D(n645), .CK(clk), .Q(dori_o) );
  DFFRHQ \decider/addrT_reg[0]  ( .D(n660), .CK(clk), .RN(rstn), .Q(addrT[0])
         );
  DFFRHQ \decider/addrT_reg[1]  ( .D(n659), .CK(clk), .RN(rstn), .Q(addrT[1])
         );
  DFFRHQ \decider/addrT_reg[2]  ( .D(n658), .CK(clk), .RN(rstn), .Q(addrT[2])
         );
  DFFRHQ \decider/addrT_reg[3]  ( .D(n657), .CK(clk), .RN(rstn), .Q(addrT[3])
         );
  DFFRHQ \decider/addrT_reg[4]  ( .D(n656), .CK(clk), .RN(rstn), .Q(addrT[4])
         );
  DFFRHQ \decider/addrT_reg[5]  ( .D(n655), .CK(clk), .RN(rstn), .Q(addrT[5])
         );
  DFFRHQ \decider/addrT_reg[6]  ( .D(n653), .CK(clk), .RN(rstn), .Q(addrT[6])
         );
  DFFRHQ \decider/addrT_reg[7]  ( .D(n652), .CK(clk), .RN(rstn), .Q(addrT[7])
         );
  DFFRHQ \decider/addrT_reg[8]  ( .D(n651), .CK(clk), .RN(rstn), .Q(addrT[8])
         );
  DFFRHQ \decider/addrT_reg[9]  ( .D(n650), .CK(clk), .RN(rstn), .Q(addrT[9])
         );
  DFFHQ \driver/db_o_reg[6]  ( .D(n377), .CK(clk), .Q(db_o[6]) );
  DFFHQ \driver/db_o_reg[5]  ( .D(n378), .CK(clk), .Q(db_o[5]) );
  DFFHQ \driver/db_o_reg[4]  ( .D(n379), .CK(clk), .Q(db_o[4]) );
  DFFHQ \driver/db_o_reg[3]  ( .D(n380), .CK(clk), .Q(db_o[3]) );
  DFFHQ \driver/db_o_reg[2]  ( .D(n646), .CK(clk), .Q(db_o[2]) );
  DFFHQ \driver/db_o_reg[1]  ( .D(n647), .CK(clk), .Q(db_o[1]) );
  DFFHQ \driver/db_o_reg[0]  ( .D(n357), .CK(clk), .Q(db_o[0]) );
  DFFHQ \driver/db_o_reg[7]  ( .D(n648), .CK(clk), .Q(db_o[7]) );
  DFFRHQ \clock_divider/cnt5k_reg[11]  ( .D(\clock_divider/N29 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[11] ) );
  DFFRHQ \clock_divider/cnt5k_reg[0]  ( .D(\clock_divider/N18 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[0] ) );
  DFFRHQ \clock_divider/cnt5k_reg[1]  ( .D(\clock_divider/N19 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[1] ) );
  DFFRHQ \clock_divider/cnt5k_reg[2]  ( .D(\clock_divider/N20 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[2] ) );
  DFFRHQ \clock_divider/cnt5k_reg[3]  ( .D(\clock_divider/N21 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[3] ) );
  DFFRHQ \clock_divider/cnt5k_reg[4]  ( .D(\clock_divider/N22 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[4] ) );
  DFFRHQ \clock_divider/cnt5k_reg[5]  ( .D(\clock_divider/N23 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[5] ) );
  DFFRHQ \clock_divider/cnt5k_reg[6]  ( .D(\clock_divider/N24 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[6] ) );
  DFFRHQ \clock_divider/cnt5k_reg[7]  ( .D(\clock_divider/N25 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[7] ) );
  DFFRHQ \clock_divider/cnt5k_reg[8]  ( .D(\clock_divider/N26 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[8] ) );
  DFFRHQ \clock_divider/cnt5k_reg[9]  ( .D(\clock_divider/N27 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[9] ) );
  DFFRHQ \clock_divider/cnt5k_reg[10]  ( .D(\clock_divider/N28 ), .CK(clk), 
        .RN(rstn), .Q(\clock_divider/cnt5k[10] ) );
  ADDF \r51/U2_1  ( .A(n669), .B(n333), .CI(\r51/carry[1] ), .CO(
        \r51/carry[2] ), .S(\decider/N88 ) );
  ADDF \r51/U2_2  ( .A(n668), .B(n332), .CI(\r51/carry[2] ), .CO(
        \r51/carry[3] ), .S(\decider/N89 ) );
  ADDF \r51/U2_3  ( .A(n667), .B(n331), .CI(\r51/carry[3] ), .CO(
        \r51/carry[4] ), .S(\decider/N90 ) );
  ADDF \r51/U2_4  ( .A(n666), .B(n330), .CI(\r51/carry[4] ), .CO(
        \r51/carry[5] ), .S(\decider/N91 ) );
  ADDF \r51/U2_5  ( .A(n665), .B(n329), .CI(\r51/carry[5] ), .CO(
        \r51/carry[6] ), .S(\decider/N92 ) );
  ADDF \r51/U2_6  ( .A(n664), .B(n654), .CI(\r51/carry[6] ), .CO(
        \r51/carry[7] ), .S(\decider/N93 ) );
  ADDF \r51/U2_7  ( .A(n663), .B(n654), .CI(\r51/carry[7] ), .CO(
        \r51/carry[8] ), .S(\decider/N94 ) );
  ADDF \r51/U2_8  ( .A(n662), .B(n654), .CI(\r51/carry[8] ), .CO(
        \r51/carry[9] ), .S(\decider/N95 ) );
  ADDF \r51/U2_9  ( .A(n661), .B(n654), .CI(\r51/carry[9] ), .S(\decider/N96 )
         );
  ADDF \r62/S3_2_3  ( .A(n673), .B(n427), .CI(n674), .CO(\r62/CARRYB[2][3] ), 
        .S(\r62/SUMB[2][3] ) );
  ADDF \r62/S2_2_2  ( .A(\r62/ab[2][2] ), .B(n426), .CI(\r62/SUMB[1][3] ), 
        .CO(\r62/CARRYB[2][2] ), .S(\r62/SUMB[2][2] ) );
  ADDF \r62/S3_3_3  ( .A(n672), .B(\r62/CARRYB[2][3] ), .CI(n673), .CO(
        \r62/CARRYB[3][3] ), .S(\r62/SUMB[3][3] ) );
  ADDF \r62/S2_3_2  ( .A(\r62/ab[3][2] ), .B(\r62/CARRYB[2][2] ), .CI(
        \r62/SUMB[2][3] ), .CO(\r62/CARRYB[3][2] ), .S(\r62/SUMB[3][2] ) );
  ADDF \r62/S1_3_0  ( .A(\r62/ab[3][0] ), .B(n425), .CI(\r62/SUMB[1][2] ), 
        .CO(\r62/CARRYB[3][0] ), .S(\decider/N58 ) );
  ADDF \r62/S3_4_3  ( .A(n671), .B(\r62/CARRYB[3][3] ), .CI(n672), .CO(
        \r62/CARRYB[4][3] ), .S(\r62/SUMB[4][3] ) );
  ADDF \r62/S2_4_2  ( .A(\r62/ab[4][2] ), .B(\r62/CARRYB[3][2] ), .CI(
        \r62/SUMB[3][3] ), .CO(\r62/CARRYB[4][2] ), .S(\r62/SUMB[4][2] ) );
  ADDF \r62/S1_4_0  ( .A(\r62/ab[4][0] ), .B(\r62/CARRYB[3][0] ), .CI(
        \r62/SUMB[2][2] ), .CO(\r62/CARRYB[4][0] ), .S(\r62/PROD1[4] ) );
  ADDF \r62/S3_5_3  ( .A(\r62/ab[7][2] ), .B(\r62/CARRYB[4][3] ), .CI(n671), 
        .CO(\r62/SUMB[6][3] ), .S(\r62/SUMB[5][3] ) );
  ADDF \r62/S2_5_2  ( .A(\r62/ab[7][2] ), .B(\r62/CARRYB[4][2] ), .CI(
        \r62/SUMB[4][3] ), .CO(\r62/CARRYB[5][2] ), .S(\r62/SUMB[5][2] ) );
  ADDF \r62/S2_6_2  ( .A(\r62/ab[7][2] ), .B(\r62/CARRYB[5][2] ), .CI(
        \r62/SUMB[5][3] ), .CO(\r62/CARRYB[6][2] ), .S(\r62/SUMB[6][2] ) );
  ADDF \r62/S2_7_2  ( .A(\r62/ab[7][2] ), .B(\r62/CARRYB[6][2] ), .CI(
        \r62/SUMB[6][3] ), .S(\r62/SUMB[7][2] ) );
  AND2 U338 ( .A(addrD[7]), .B(addrD[6]), .Y(n401) );
  AND2 U339 ( .A(addrD[8]), .B(n401), .Y(n402) );
  AND2 U340 ( .A(\clock_divider/cnt5k[10] ), .B(n410), .Y(n403) );
  AND2 U341 ( .A(\clock_divider/cnt5k[8] ), .B(n411), .Y(n404) );
  AND2 U342 ( .A(\clock_divider/cnt5k[6] ), .B(n412), .Y(n405) );
  AND2 U343 ( .A(\clock_divider/cnt5k[4] ), .B(n413), .Y(n406) );
  AND2 U344 ( .A(\clock_divider/cnt5k[2] ), .B(n414), .Y(n407) );
  AND2 U345 ( .A(\add_2_root_decider/add_109_3_cf/carry[4] ), .B(
        \r62/PROD1[4] ), .Y(n408) );
  AND2 U346 ( .A(n682), .B(\sub_1_root_decider/sub_49/carry[3] ), .Y(n409) );
  AND2 U347 ( .A(\clock_divider/cnt5k[9] ), .B(n404), .Y(n410) );
  AND2 U348 ( .A(\clock_divider/cnt5k[7] ), .B(n405), .Y(n411) );
  AND2 U349 ( .A(\clock_divider/cnt5k[5] ), .B(n406), .Y(n412) );
  AND2 U350 ( .A(\clock_divider/cnt5k[3] ), .B(n407), .Y(n413) );
  AND2 U351 ( .A(\clock_divider/cnt5k[1] ), .B(\clock_divider/cnt5k[0] ), .Y(
        n414) );
  AND2 U352 ( .A(\add_2_root_decider/add_109_3_cf/carry[7] ), .B(\decider/N62 ), .Y(n415) );
  AND2 U353 ( .A(n682), .B(n681), .Y(n416) );
  AND2 U354 ( .A(\r62/CARRYB[4][0] ), .B(\r62/SUMB[3][2] ), .Y(n417) );
  AND2 U355 ( .A(n417), .B(\r62/SUMB[4][2] ), .Y(n418) );
  AND2 U356 ( .A(n418), .B(\r62/SUMB[5][2] ), .Y(n419) );
  OR2 U357 ( .A(n626), .B(n562), .Y(n420) );
  AND2 U358 ( .A(addrD[9]), .B(n402), .Y(n421) );
  AND2 U359 ( .A(\clock_divider/cnt5k[11] ), .B(n403), .Y(n422) );
  AND2 U360 ( .A(n415), .B(\decider/N63 ), .Y(n423) );
  AND2 U361 ( .A(n419), .B(\r62/SUMB[6][2] ), .Y(n424) );
  AND2 U362 ( .A(\r62/ab[2][0] ), .B(\r62/ab[0][2] ), .Y(n425) );
  AND2 U363 ( .A(n675), .B(\r62/ab[1][2] ), .Y(n426) );
  AND2 U364 ( .A(n675), .B(n674), .Y(n427) );
  BUF U365 ( .I(n545), .O(n428) );
  INV U366 ( .A(n463), .Y(n429) );
  INV U367 ( .A(n576), .Y(n430) );
  BUF U368 ( .I(n521), .O(n431) );
  BUF U369 ( .I(n466), .O(n432) );
  BUF U370 ( .I(n635), .O(n433) );
  BUF U371 ( .I(n456), .O(n434) );
  BUF U372 ( .I(n456), .O(n435) );
  LOGIC_0 U373 ( .LOGIC_0_PIN(\driver/*Logic0* ) );
  NAND2 U374 ( .A(n436), .B(n437), .Y(\r51/carry[1] ) );
  XNOR2 U375 ( .A(n334), .B(n670), .Y(\decider/N38 ) );
  INV U376 ( .A(n334), .Y(n436) );
  INV U377 ( .A(n670), .Y(n437) );
  NAND2 U378 ( .A(n438), .B(n439), .Y(
        \add_2_root_decider/add_109_3_cf/carry[2] ) );
  XNOR2 U379 ( .A(\r62/ab[1][0] ), .B(\decider/N55 ), .Y(\decider/N85 ) );
  INV U380 ( .A(\r62/ab[1][0] ), .Y(n438) );
  INV U381 ( .A(\decider/N55 ), .Y(n439) );
  NAND2 U382 ( .A(n440), .B(n449), .Y(
        \add_2_root_decider/add_109_3_cf/carry[4] ) );
  XNOR2 U383 ( .A(\decider/N58 ), .B(
        \add_2_root_decider/add_109_3_cf/carry[3] ), .Y(\decider/N83 ) );
  INV U384 ( .A(\decider/N58 ), .Y(n440) );
  NAND2 U385 ( .A(n441), .B(n450), .Y(
        \add_2_root_decider/add_109_3_cf/carry[7] ) );
  XNOR2 U386 ( .A(\decider/N61 ), .B(
        \add_2_root_decider/add_109_3_cf/carry[6] ), .Y(\decider/N80 ) );
  INV U387 ( .A(\decider/N61 ), .Y(n441) );
  NAND2 U388 ( .A(addrD[1]), .B(addrD[0]), .Y(
        \sub_1_root_decider/sub_49/carry[2] ) );
  XNOR2 U389 ( .A(n680), .B(n679), .Y(\decider/posy_m_rex_top[1] ) );
  NAND2 U390 ( .A(addrD[2]), .B(n442), .Y(\sub_1_root_decider/sub_49/carry[3] ) );
  XNOR2 U391 ( .A(n681), .B(\sub_1_root_decider/sub_49/carry[2] ), .Y(
        \decider/posy_m_rex_top[2] ) );
  INV U392 ( .A(\sub_1_root_decider/sub_49/carry[2] ), .Y(n442) );
  NAND2 U393 ( .A(addrD[5]), .B(n451), .Y(\sub_1_root_decider/sub_49/carry[6] ) );
  XNOR2 U394 ( .A(n678), .B(\sub_1_root_decider/sub_49/carry[5] ), .Y(
        \decider/posy_m_rex_top[5] ) );
  NAND2 U395 ( .A(n544), .B(n443), .Y(\decider/sub_45/carry[5] ) );
  XNOR2 U396 ( .A(addrD[10]), .B(\decider/sub_45/carry[4] ), .Y(
        \decider/posx_m_rex_left [7]) );
  INV U397 ( .A(\decider/sub_45/carry[4] ), .Y(n443) );
  NAND2 U398 ( .A(n444), .B(n445), .Y(\decider/sub_45/carry[4] ) );
  XNOR2 U399 ( .A(addrD[9]), .B(\decider/sub_45/carry[3] ), .Y(
        \decider/posx_m_rex_left [6]) );
  INV U400 ( .A(addrD[9]), .Y(n444) );
  INV U401 ( .A(\decider/sub_45/carry[3] ), .Y(n445) );
  NAND2 U402 ( .A(n547), .B(n446), .Y(\decider/sub_45/carry[3] ) );
  XNOR2 U403 ( .A(addrD[8]), .B(\decider/sub_45/carry[2] ), .Y(
        \decider/posx_m_rex_left [5]) );
  INV U404 ( .A(\decider/sub_45/carry[2] ), .Y(n446) );
  NAND2 U405 ( .A(n447), .B(n675), .Y(\decider/sub_45/carry[2] ) );
  XNOR2 U406 ( .A(addrD[7]), .B(addrD[6]), .Y(\decider/posx_m_rex_left [4]) );
  INV U407 ( .A(addrD[7]), .Y(n447) );
  NAND2 U408 ( .A(addrD[5]), .B(n452), .Y(\decider/sub_75/carry[6] ) );
  XNOR2 U409 ( .A(n678), .B(\decider/sub_75/carry[5] ), .Y(
        \decider/posy_m_obstacle_top [5]) );
  XNOR2 U410 ( .A(n677), .B(\sub_0_root_decider/sub_73/carry[15] ), .Y(
        \decider/posx_m_obstacle_right[15] ) );
  NAND2 U411 ( .A(n444), .B(n453), .Y(\r187/carry[7] ) );
  XNOR2 U412 ( .A(addrD[9]), .B(n402), .Y(\decider/obstacle_right [6]) );
  NAND2 U413 ( .A(n544), .B(n448), .Y(\r187/carry[8] ) );
  XNOR2 U414 ( .A(addrD[10]), .B(\r187/carry[7] ), .Y(
        \decider/obstacle_right [7]) );
  INV U415 ( .A(\r187/carry[7] ), .Y(n448) );
  XOR2 U416 ( .A(addrD[7]), .B(addrD[6]), .Y(\driver/N44 ) );
  XOR2 U417 ( .A(addrD[8]), .B(n401), .Y(\driver/N45 ) );
  XOR2 U418 ( .A(addrD[9]), .B(n402), .Y(\driver/N46 ) );
  XOR2 U419 ( .A(addrD[10]), .B(n421), .Y(\driver/N47 ) );
  XOR2 U420 ( .A(\clock_divider/cnt5k[12] ), .B(n422), .Y(\clock_divider/N17 )
         );
  XOR2 U421 ( .A(\clock_divider/cnt5k[11] ), .B(n403), .Y(\clock_divider/N16 )
         );
  XOR2 U422 ( .A(\clock_divider/cnt5k[10] ), .B(n410), .Y(\clock_divider/N15 )
         );
  XOR2 U423 ( .A(\clock_divider/cnt5k[9] ), .B(n404), .Y(\clock_divider/N14 )
         );
  XOR2 U424 ( .A(\clock_divider/cnt5k[8] ), .B(n411), .Y(\clock_divider/N13 )
         );
  XOR2 U425 ( .A(\clock_divider/cnt5k[7] ), .B(n405), .Y(\clock_divider/N12 )
         );
  XOR2 U426 ( .A(\clock_divider/cnt5k[6] ), .B(n412), .Y(\clock_divider/N11 )
         );
  XOR2 U427 ( .A(\clock_divider/cnt5k[5] ), .B(n406), .Y(\clock_divider/N10 )
         );
  XOR2 U428 ( .A(\clock_divider/cnt5k[4] ), .B(n413), .Y(\clock_divider/N9 )
         );
  XOR2 U429 ( .A(\clock_divider/cnt5k[3] ), .B(n407), .Y(\clock_divider/N8 )
         );
  XOR2 U430 ( .A(\clock_divider/cnt5k[2] ), .B(n414), .Y(\clock_divider/N7 )
         );
  XOR2 U431 ( .A(\clock_divider/cnt5k[1] ), .B(\clock_divider/cnt5k[0] ), .Y(
        \clock_divider/N6 ) );
  XOR2 U432 ( .A(\decider/N57 ), .B(\add_2_root_decider/add_109_3_cf/carry[2] ), .Y(\decider/N84 ) );
  NAND2 U433 ( .A(\add_2_root_decider/add_109_3_cf/carry[2] ), .B(
        \decider/N57 ), .Y(n449) );
  INV U434 ( .A(n449), .Y(\add_2_root_decider/add_109_3_cf/carry[3] ) );
  XOR2 U435 ( .A(\r62/PROD1[4] ), .B(
        \add_2_root_decider/add_109_3_cf/carry[4] ), .Y(\decider/N82 ) );
  XOR2 U436 ( .A(\decider/N60 ), .B(n408), .Y(\decider/N81 ) );
  NAND2 U437 ( .A(n408), .B(\decider/N60 ), .Y(n450) );
  INV U438 ( .A(n450), .Y(\add_2_root_decider/add_109_3_cf/carry[6] ) );
  XOR2 U439 ( .A(\decider/N62 ), .B(\add_2_root_decider/add_109_3_cf/carry[7] ), .Y(\decider/N79 ) );
  XOR2 U440 ( .A(\decider/N63 ), .B(n415), .Y(\decider/N78 ) );
  XOR2 U441 ( .A(\decider/N64 ), .B(n423), .Y(\decider/N77 ) );
  XOR2 U442 ( .A(\r62/ab[1][2] ), .B(n675), .Y(\r62/SUMB[1][2] ) );
  XOR2 U443 ( .A(n674), .B(n675), .Y(\r62/SUMB[1][3] ) );
  XOR2 U444 ( .A(n682), .B(\sub_1_root_decider/sub_49/carry[3] ), .Y(
        \decider/posy_m_rex_top[3] ) );
  XOR2 U445 ( .A(n676), .B(n409), .Y(\decider/posy_m_rex_top[4] ) );
  NAND2 U446 ( .A(n676), .B(n409), .Y(n451) );
  INV U447 ( .A(n451), .Y(\sub_1_root_decider/sub_49/carry[5] ) );
  XOR2 U448 ( .A(n682), .B(n681), .Y(\decider/posy_m_obstacle_top [3]) );
  XOR2 U449 ( .A(n676), .B(n416), .Y(\decider/posy_m_obstacle_top [4]) );
  NAND2 U450 ( .A(n676), .B(n416), .Y(n452) );
  INV U451 ( .A(n452), .Y(\decider/sub_75/carry[5] ) );
  XOR2 U452 ( .A(addrD[8]), .B(n401), .Y(\decider/obstacle_right [5]) );
  NAND2 U453 ( .A(addrD[8]), .B(n401), .Y(n453) );
  XOR2 U454 ( .A(\r62/ab[2][0] ), .B(\r62/ab[0][2] ), .Y(\decider/N57 ) );
  XOR2 U455 ( .A(\r62/CARRYB[4][0] ), .B(\r62/SUMB[3][2] ), .Y(\decider/N60 )
         );
  XOR2 U456 ( .A(n417), .B(\r62/SUMB[4][2] ), .Y(\decider/N61 ) );
  XOR2 U457 ( .A(n418), .B(\r62/SUMB[5][2] ), .Y(\decider/N62 ) );
  XOR2 U458 ( .A(n419), .B(\r62/SUMB[6][2] ), .Y(\decider/N63 ) );
  XOR2 U459 ( .A(n424), .B(\r62/SUMB[7][2] ), .Y(\decider/N64 ) );
  INV U460 ( .A(n454), .Y(\sub_0_root_decider/sub_73/carry[15] ) );
  NOR4BB U461 ( .AN(n455), .BN(\r187/carry[8] ), .C(
        \decider/obstacle_right [5]), .D(\driver/N44 ), .Y(n454) );
  NOR2 U462 ( .A(\decider/obstacle_right [7]), .B(\decider/obstacle_right [6]), 
        .Y(n455) );
  NOR2B U463 ( .AN(n671), .B(n435), .Y(\r62/ab[4][2] ) );
  NOR2B U464 ( .AN(n671), .B(n457), .Y(\r62/ab[4][0] ) );
  NOR2B U465 ( .AN(n672), .B(n434), .Y(\r62/ab[3][2] ) );
  NOR2B U466 ( .AN(n672), .B(n457), .Y(\r62/ab[3][0] ) );
  NOR2B U467 ( .AN(n673), .B(n435), .Y(\r62/ab[2][2] ) );
  NOR2B U468 ( .AN(n673), .B(n457), .Y(\r62/ab[2][0] ) );
  NOR2B U469 ( .AN(n674), .B(n434), .Y(\r62/ab[1][2] ) );
  NOR2B U470 ( .AN(n675), .B(n435), .Y(\r62/ab[0][2] ) );
  OAI2BB1 U471 ( .A0N(n458), .A1N(dori_o), .B0(n459), .Y(n645) );
  NOR2B U472 ( .AN(n460), .B(n461), .Y(n458) );
  OAI211 U473 ( .A0(n462), .A1(n463), .B0(n464), .C0(n465), .Y(n646) );
  AOI222 U474 ( .A0(db_o[2]), .A1(n432), .B0(addrD[8]), .B1(n467), .C0(n468), 
        .C1(addrD[2]), .Y(n465) );
  AOI2BB1 U475 ( .A0N(n469), .A1N(n470), .B0(n471), .Y(n464) );
  AOI32 U476 ( .A0(n472), .A1(n473), .A2(n474), .B0(n475), .B1(addrT[1]), .Y(
        n469) );
  AOI211 U477 ( .A0(n476), .A1(n477), .B0(n478), .C0(n479), .Y(n462) );
  OAI2BB1 U478 ( .A0N(n480), .A1N(n481), .B0(n482), .Y(n476) );
  OAI211 U479 ( .A0(n483), .A1(n463), .B0(n484), .C0(n485), .Y(n647) );
  AOI222 U480 ( .A0(db_o[1]), .A1(n432), .B0(addrD[7]), .B1(n467), .C0(n468), 
        .C1(addrD[1]), .Y(n485) );
  AOI31 U481 ( .A0(n486), .A1(n473), .A2(n487), .B0(n471), .Y(n484) );
  NOR2B U482 ( .AN(n474), .B(n470), .Y(n487) );
  NOR4 U483 ( .A(n488), .B(n489), .C(n490), .D(n491), .Y(n483) );
  OAI2BB2 U484 ( .B0(n492), .B1(n493), .A0N(n494), .A1N(n495), .Y(n491) );
  OAI32 U485 ( .A0(n496), .A1(addrT[3]), .A2(n497), .B0(n498), .B1(n499), .Y(
        n489) );
  AOI21 U486 ( .A0(addrT[4]), .A1(n500), .B0(n501), .Y(n498) );
  OAI21 U487 ( .A0(addrT[0]), .A1(n502), .B0(n503), .Y(n500) );
  OAI31 U488 ( .A0(n504), .A1(n505), .A2(n506), .B0(n507), .Y(n488) );
  INV U489 ( .A(n508), .Y(n507) );
  INV U490 ( .A(n509), .Y(n648) );
  AOI221 U491 ( .A0(n510), .A1(n511), .B0(n432), .B1(db_o[7]), .C0(n467), .Y(
        n509) );
  OAI211 U492 ( .A0(n496), .A1(n512), .B0(n513), .C0(n514), .Y(n510) );
  AOI31 U493 ( .A0(n515), .A1(n502), .A2(n486), .B0(n516), .Y(n513) );
  INV U494 ( .A(n517), .Y(n516) );
  OAI31 U495 ( .A0(n518), .A1(n519), .A2(n481), .B0(n480), .Y(n517) );
  MX2 U496 ( .A(addrT[3]), .B(addrT[4]), .S0(n430), .Y(n518) );
  MX2 U497 ( .A(\decider/N96 ), .B(addrT[9]), .S0(n431), .Y(n650) );
  MX2 U498 ( .A(\decider/N95 ), .B(addrT[8]), .S0(n431), .Y(n651) );
  MX2 U499 ( .A(\decider/N94 ), .B(addrT[7]), .S0(n431), .Y(n652) );
  MX2 U500 ( .A(\decider/N93 ), .B(addrT[6]), .S0(n431), .Y(n653) );
  NOR2B U501 ( .AN(\decider/sub_75/carry[6] ), .B(n434), .Y(n654) );
  MX2 U502 ( .A(\decider/N92 ), .B(addrT[5]), .S0(n431), .Y(n655) );
  MX2 U503 ( .A(\decider/N91 ), .B(addrT[4]), .S0(n431), .Y(n656) );
  MX2 U504 ( .A(\decider/N90 ), .B(addrT[3]), .S0(n431), .Y(n657) );
  MX2 U505 ( .A(\decider/N89 ), .B(addrT[2]), .S0(n431), .Y(n658) );
  MX2 U506 ( .A(\decider/N88 ), .B(addrT[1]), .S0(n431), .Y(n659) );
  MX2 U507 ( .A(\decider/N38 ), .B(addrT[0]), .S0(n431), .Y(n660) );
  AOI31 U508 ( .A0(\decider/posx_m_obstacle_right[15] ), .A1(n522), .A2(
        \r187/carry[8] ), .B0(n435), .Y(n521) );
  INV U509 ( .A(\decider/sub_75/carry[6] ), .Y(n522) );
  MX2 U510 ( .A(\decider/N77 ), .B(\decider/N64 ), .S0(n435), .Y(n661) );
  MX2 U511 ( .A(\decider/N78 ), .B(\decider/N63 ), .S0(n434), .Y(n662) );
  MX2 U512 ( .A(\decider/N79 ), .B(\decider/N62 ), .S0(n435), .Y(n663) );
  MX2 U513 ( .A(\decider/N80 ), .B(\decider/N61 ), .S0(n434), .Y(n664) );
  MX2 U514 ( .A(\decider/N81 ), .B(\decider/N60 ), .S0(n435), .Y(n665) );
  MX2 U515 ( .A(\decider/N82 ), .B(\r62/PROD1[4] ), .S0(n434), .Y(n666) );
  MX2 U516 ( .A(\decider/N83 ), .B(\decider/N58 ), .S0(n435), .Y(n667) );
  MX2 U517 ( .A(\decider/N84 ), .B(\decider/N57 ), .S0(n434), .Y(n668) );
  OAI2BB1 U518 ( .A0N(\decider/N85 ), .A1N(n457), .B0(n438), .Y(n669) );
  NOR2B U519 ( .AN(n674), .B(n457), .Y(\r62/ab[1][0] ) );
  INV U520 ( .A(n434), .Y(n457) );
  NAND2 U521 ( .A(n435), .B(addrD[6]), .Y(n670) );
  MX2 U522 ( .A(\decider/obstacle_right [7]), .B(\decider/posx_m_rex_left [7]), 
        .S0(n435), .Y(n671) );
  MX2 U523 ( .A(\decider/obstacle_right [6]), .B(\decider/posx_m_rex_left [6]), 
        .S0(n434), .Y(n672) );
  MX2 U524 ( .A(\decider/obstacle_right [5]), .B(\decider/posx_m_rex_left [5]), 
        .S0(n435), .Y(n673) );
  MX2 U525 ( .A(\driver/N44 ), .B(\decider/posx_m_rex_left [4]), .S0(n434), 
        .Y(n674) );
  INV U526 ( .A(addrD[4]), .Y(n676) );
  MX2 U527 ( .A(n523), .B(n524), .S0(addrD[5]), .Y(n397) );
  OAI21 U528 ( .A0(addrD[4]), .A1(n459), .B0(n525), .Y(n524) );
  NOR2 U529 ( .A(n459), .B(n526), .Y(n523) );
  MX2 U530 ( .A(n527), .B(n460), .S0(addrD[0]), .Y(n396) );
  MX2 U531 ( .A(n528), .B(n529), .S0(addrD[1]), .Y(n395) );
  INV U532 ( .A(n530), .Y(n529) );
  NOR2B U533 ( .AN(addrD[0]), .B(n459), .Y(n528) );
  MX2 U534 ( .A(n531), .B(n532), .S0(addrD[2]), .Y(n394) );
  OAI21 U535 ( .A0(addrD[1]), .A1(n459), .B0(n530), .Y(n532) );
  AOI2BB1 U536 ( .A0N(addrD[0]), .A1N(n459), .B0(n460), .Y(n530) );
  NOR3B U537 ( .AN(addrD[1]), .B(n459), .C(n679), .Y(n531) );
  MX2 U538 ( .A(n533), .B(n534), .S0(addrD[3]), .Y(n393) );
  NOR2B U539 ( .AN(n535), .B(n459), .Y(n533) );
  MX2 U540 ( .A(n536), .B(n537), .S0(addrD[4]), .Y(n392) );
  INV U541 ( .A(n525), .Y(n537) );
  AOI2BB1 U542 ( .A0N(addrD[3]), .A1N(n459), .B0(n534), .Y(n525) );
  OAI21 U543 ( .A0(n535), .A1(n459), .B0(n538), .Y(n534) );
  NOR3B U544 ( .AN(n535), .B(n459), .C(n682), .Y(n536) );
  INV U545 ( .A(addrD[3]), .Y(n682) );
  INV U546 ( .A(n527), .Y(n459) );
  NOR3B U547 ( .AN(n539), .B(n460), .C(n649), .Y(n527) );
  INV U548 ( .A(n538), .Y(n460) );
  OAI21 U549 ( .A0(n540), .A1(n541), .B0(n542), .Y(n538) );
  OAI2BB2 U550 ( .B0(n543), .B1(n544), .A0N(\driver/N47 ), .A1N(n428), .Y(n391) );
  MX2 U551 ( .A(n428), .B(n546), .S0(addrD[6]), .Y(n390) );
  OAI2BB2 U552 ( .B0(n447), .B1(n543), .A0N(\driver/N44 ), .A1N(n428), .Y(n389) );
  OAI2BB2 U553 ( .B0(n547), .B1(n543), .A0N(\driver/N45 ), .A1N(n428), .Y(n388) );
  OAI2BB2 U554 ( .B0(n543), .B1(n444), .A0N(\driver/N46 ), .A1N(n428), .Y(n387) );
  NOR3B U555 ( .AN(rstn), .B(n546), .C(n548), .Y(n545) );
  INV U556 ( .A(n543), .Y(n546) );
  OAI21 U557 ( .A0(n549), .A1(n550), .B0(n551), .Y(n386) );
  NAND2 U558 ( .A(n552), .B(n551), .Y(n385) );
  MX2 U559 ( .A(n553), .B(n554), .S0(n555), .Y(n552) );
  AOI31 U560 ( .A0(cs_o[3]), .A1(addrD[7]), .A2(n556), .B0(n557), .Y(n553) );
  NOR3B U561 ( .AN(addrD[6]), .B(n547), .C(n548), .Y(n556) );
  INV U562 ( .A(addrD[8]), .Y(n547) );
  NAND3B U563 ( .AN(n558), .B(n551), .C(n559), .Y(n384) );
  MX2 U564 ( .A(n548), .B(n560), .S0(n555), .Y(n559) );
  OAI31 U565 ( .A0(n561), .A1(n649), .A2(n562), .B0(n550), .Y(n551) );
  INV U566 ( .A(n555), .Y(n550) );
  AOI211 U567 ( .A0(en_o), .A1(n561), .B0(n461), .C0(n543), .Y(n555) );
  OAI32 U568 ( .A0(n542), .A1(n678), .A2(n526), .B0(n541), .B1(n540), .Y(n543)
         );
  NOR2 U569 ( .A(n649), .B(n563), .Y(n540) );
  NOR2B U570 ( .AN(\driver/start_history [1]), .B(start), .Y(n563) );
  NAND3 U571 ( .A(addrD[4]), .B(n535), .C(addrD[3]), .Y(n526) );
  NOR3B U572 ( .AN(addrD[1]), .B(n679), .C(n681), .Y(n535) );
  INV U573 ( .A(addrD[2]), .Y(n681) );
  INV U574 ( .A(addrD[0]), .Y(n679) );
  INV U575 ( .A(addrD[5]), .Y(n678) );
  INV U576 ( .A(n564), .Y(n542) );
  NOR2B U577 ( .AN(state[2]), .B(n558), .Y(n561) );
  INV U578 ( .A(n565), .Y(n380) );
  AOI221 U579 ( .A0(n468), .A1(addrD[3]), .B0(db_o[3]), .B1(n432), .C0(n566), 
        .Y(n565) );
  OAI221 U580 ( .A0(n567), .A1(n470), .B0(n568), .B1(n463), .C0(n569), .Y(n566) );
  NOR4BB U581 ( .AN(n570), .BN(n482), .C(n571), .D(n572), .Y(n568) );
  NOR3B U582 ( .AN(n477), .B(n496), .C(n573), .Y(n572) );
  AOI221 U583 ( .A0(n574), .A1(n575), .B0(n576), .B1(n479), .C0(n478), .Y(n570) );
  OAI221 U584 ( .A0(n577), .A1(n578), .B0(n496), .B1(n493), .C0(n579), .Y(n478) );
  AOI2BB2 U585 ( .B0(n506), .B1(n503), .A0N(n473), .A1N(n520), .Y(n577) );
  AOI22 U586 ( .A0(n497), .A1(n580), .B0(n475), .B1(n520), .Y(n567) );
  INV U587 ( .A(n581), .Y(n379) );
  AOI221 U588 ( .A0(n468), .A1(addrD[4]), .B0(db_o[4]), .B1(n432), .C0(n582), 
        .Y(n581) );
  OAI221 U589 ( .A0(n583), .A1(n470), .B0(n584), .B1(n463), .C0(n569), .Y(n582) );
  NOR4B U590 ( .AN(n579), .B(n571), .C(n585), .D(n586), .Y(n584) );
  OAI32 U591 ( .A0(n492), .A1(addrT[5]), .A2(n587), .B0(n588), .B1(n482), .Y(
        n586) );
  AOI2BB1 U592 ( .A0N(addrT[3]), .A1N(n502), .B0(n519), .Y(n588) );
  AOI2BB2 U593 ( .B0(addrT[4]), .B1(n589), .A0N(n576), .A1N(n493), .Y(n587) );
  OAI2BB1 U594 ( .A0N(addrT[2]), .A1N(n576), .B0(n504), .Y(n589) );
  AOI2BB1 U595 ( .A0N(n590), .A1N(n479), .B0(addrT[1]), .Y(n585) );
  NOR2 U596 ( .A(n508), .B(n591), .Y(n579) );
  AOI2BB2 U597 ( .B0(n494), .B1(n502), .A0N(n477), .A1N(n592), .Y(n583) );
  OAI211 U598 ( .A0(n593), .A1(n463), .B0(n569), .C0(n594), .Y(n378) );
  AOI22 U599 ( .A0(db_o[5]), .A1(n432), .B0(addrD[5]), .B1(n468), .Y(n594) );
  NAND2 U600 ( .A(n420), .B(n595), .Y(n569) );
  NOR2B U601 ( .AN(n596), .B(n597), .Y(n593) );
  OAI221 U602 ( .A0(n598), .A1(n512), .B0(n482), .B1(n504), .C0(n599), .Y(n597) );
  AOI221 U603 ( .A0(n600), .A1(n520), .B0(n494), .B1(n575), .C0(n601), .Y(n598) );
  OAI221 U604 ( .A0(n602), .A1(n496), .B0(n492), .B1(n573), .C0(n603), .Y(n601) );
  OR4 U605 ( .A(n604), .B(n502), .C(n473), .D(addrT[0]), .Y(n603) );
  INV U606 ( .A(n486), .Y(n492) );
  NOR2B U607 ( .AN(n477), .B(n506), .Y(n602) );
  AOI211 U608 ( .A0(n479), .A1(n575), .B0(n571), .C0(n605), .Y(n596) );
  NOR4BB U609 ( .AN(addrT[0]), .BN(addrT[2]), .C(n604), .D(n573), .Y(n605) );
  NAND2B U610 ( .AN(n473), .B(n502), .Y(n573) );
  NOR3B U611 ( .AN(n606), .B(n504), .C(addrT[0]), .Y(n571) );
  AND2 U612 ( .A(n475), .B(n607), .Y(n479) );
  NOR3B U613 ( .AN(addrT[4]), .B(n499), .C(addrT[6]), .Y(n475) );
  INV U614 ( .A(n608), .Y(n377) );
  AOI211 U615 ( .A0(n609), .A1(n511), .B0(n468), .C0(n610), .Y(n608) );
  OAI2BB2 U616 ( .B0(n470), .B1(n611), .A0N(db_o[6]), .A1N(n432), .Y(n610) );
  AOI221 U617 ( .A0(n486), .A1(n481), .B0(n506), .B1(n600), .C0(n612), .Y(n611) );
  OAI221 U618 ( .A0(n613), .A1(n474), .B0(n614), .B1(n604), .C0(n496), .Y(n612) );
  INV U619 ( .A(n472), .Y(n496) );
  NAND2 U620 ( .A(n502), .B(addrT[0]), .Y(n614) );
  NOR2B U621 ( .AN(addrT[4]), .B(n506), .Y(n481) );
  NAND2 U622 ( .A(n429), .B(addrT[3]), .Y(n470) );
  OAI31 U623 ( .A0(n604), .A1(addrT[0]), .A2(n504), .B0(n599), .Y(n609) );
  NOR4 U624 ( .A(n591), .B(n590), .C(n615), .D(n616), .Y(n599) );
  OAI31 U625 ( .A0(n592), .A1(n512), .A2(n477), .B0(n514), .Y(n616) );
  AOI211 U626 ( .A0(n472), .A1(addrT[4]), .B0(n617), .C0(n508), .Y(n514) );
  NOR2B U627 ( .AN(n574), .B(n477), .Y(n508) );
  NOR4BB U628 ( .AN(addrT[7]), .BN(n515), .C(addrT[6]), .D(n520), .Y(n617) );
  NOR3B U629 ( .AN(n607), .B(addrT[4]), .C(addrT[5]), .Y(n515) );
  NOR2B U630 ( .AN(n477), .B(addrT[3]), .Y(n607) );
  NOR2B U631 ( .AN(n486), .B(n618), .Y(n472) );
  INV U632 ( .A(n600), .Y(n592) );
  NOR3B U633 ( .AN(n473), .B(n499), .C(addrT[6]), .Y(n600) );
  INV U634 ( .A(n619), .Y(n499) );
  NOR3B U635 ( .AN(n486), .B(n493), .C(n495), .Y(n615) );
  NOR2B U636 ( .AN(n477), .B(n520), .Y(n495) );
  NOR3B U637 ( .AN(n486), .B(n473), .C(n504), .Y(n590) );
  NOR2B U638 ( .AN(addrT[6]), .B(addrT[7]), .Y(n486) );
  NOR2B U639 ( .AN(n574), .B(n576), .Y(n591) );
  NOR2B U640 ( .AN(n512), .B(n505), .Y(n574) );
  INV U641 ( .A(n606), .Y(n505) );
  INV U642 ( .A(n519), .Y(n504) );
  NOR2B U643 ( .AN(n477), .B(n512), .Y(n519) );
  INV U644 ( .A(addrT[2]), .Y(n477) );
  INV U645 ( .A(n480), .Y(n604) );
  INV U646 ( .A(n620), .Y(n357) );
  AOI221 U647 ( .A0(n468), .A1(addrD[0]), .B0(db_o[0]), .B1(n432), .C0(n621), 
        .Y(n620) );
  OAI221 U648 ( .A0(n622), .A1(n463), .B0(n675), .B1(n623), .C0(n624), .Y(n621) );
  INV U649 ( .A(n471), .Y(n624) );
  NOR2B U650 ( .AN(n562), .B(n625), .Y(n471) );
  INV U651 ( .A(n467), .Y(n623) );
  NOR2B U652 ( .AN(n626), .B(n625), .Y(n467) );
  INV U653 ( .A(addrD[6]), .Y(n675) );
  INV U654 ( .A(n511), .Y(n463) );
  NOR4 U655 ( .A(addrT[9]), .B(addrT[8]), .C(\r62/ab[7][2] ), .D(n627), .Y(
        n511) );
  OAI211 U656 ( .A0(n434), .A1(n628), .B0(n539), .C0(n595), .Y(n627) );
  NOR2B U657 ( .AN(\decider/posx_m_obstacle_right[15] ), .B(
        \decider/sub_75/carry[6] ), .Y(n628) );
  AOI211 U658 ( .A0(n619), .A1(n629), .B0(n630), .C0(n490), .Y(n622) );
  OAI21 U659 ( .A0(addrT[3]), .A1(n482), .B0(n578), .Y(n490) );
  NAND3 U660 ( .A(addrT[3]), .B(addrT[2]), .C(n619), .Y(n578) );
  OAI33 U661 ( .A0(n482), .A1(addrT[2]), .A2(n506), .B0(n613), .B1(addrT[3]), 
        .B2(n497), .Y(n630) );
  NOR2B U662 ( .AN(addrT[2]), .B(n576), .Y(n497) );
  INV U663 ( .A(n580), .Y(n613) );
  NOR2B U664 ( .AN(n480), .B(addrT[4]), .Y(n580) );
  INV U665 ( .A(n575), .Y(n506) );
  NOR2B U666 ( .AN(n502), .B(addrT[0]), .Y(n575) );
  INV U667 ( .A(n494), .Y(n482) );
  NOR2B U668 ( .AN(n606), .B(addrT[4]), .Y(n494) );
  NOR2B U669 ( .AN(n480), .B(addrT[6]), .Y(n606) );
  NOR2B U670 ( .AN(addrT[5]), .B(addrT[7]), .Y(n480) );
  OAI222 U671 ( .A0(n631), .A1(n493), .B0(n576), .B1(n632), .C0(n633), .C1(
        n473), .Y(n629) );
  AOI21 U672 ( .A0(addrT[1]), .A1(addrT[3]), .B0(addrT[6]), .Y(n633) );
  NAND2 U673 ( .A(n503), .B(addrT[3]), .Y(n632) );
  INV U674 ( .A(addrT[6]), .Y(n503) );
  INV U675 ( .A(n520), .Y(n576) );
  NOR2B U676 ( .AN(addrT[0]), .B(n502), .Y(n520) );
  INV U677 ( .A(n501), .Y(n493) );
  NOR2B U678 ( .AN(n512), .B(n473), .Y(n501) );
  INV U679 ( .A(addrT[4]), .Y(n473) );
  INV U680 ( .A(addrT[3]), .Y(n512) );
  NOR2B U681 ( .AN(n474), .B(addrT[0]), .Y(n631) );
  NOR2B U682 ( .AN(addrT[2]), .B(n502), .Y(n474) );
  INV U683 ( .A(addrT[1]), .Y(n502) );
  NOR2B U684 ( .AN(n618), .B(addrT[7]), .Y(n619) );
  INV U685 ( .A(addrT[5]), .Y(n618) );
  NOR2B U686 ( .AN(n557), .B(n625), .Y(n468) );
  INV U687 ( .A(n595), .Y(n625) );
  NOR2B U688 ( .AN(rstn), .B(n432), .Y(n595) );
  NOR3B U689 ( .AN(n541), .B(n461), .C(n564), .Y(n466) );
  NOR2B U690 ( .AN(en_o), .B(n548), .Y(n564) );
  INV U691 ( .A(n539), .Y(n548) );
  NOR3B U692 ( .AN(n554), .B(state[2]), .C(state[1]), .Y(n539) );
  AOI2BB1 U693 ( .A0N(n557), .A1N(n420), .B0(n634), .Y(n461) );
  INV U694 ( .A(en_o), .Y(n634) );
  NOR2B U695 ( .AN(n558), .B(state[2]), .Y(n562) );
  NOR3B U696 ( .AN(n549), .B(state[1]), .C(n554), .Y(n626) );
  INV U697 ( .A(state[0]), .Y(n554) );
  AOI31 U698 ( .A0(state[2]), .A1(en_o), .A2(n558), .B0(n649), .Y(n541) );
  INV U699 ( .A(rstn), .Y(n649) );
  NOR2B U700 ( .AN(state[0]), .B(n560), .Y(n558) );
  NOR3B U701 ( .AN(n549), .B(n560), .C(state[0]), .Y(n557) );
  INV U702 ( .A(state[1]), .Y(n560) );
  INV U703 ( .A(state[2]), .Y(n549) );
  XOR2 U704 ( .A(n433), .B(start), .Y(n356) );
  XOR2 U705 ( .A(addrD[0]), .B(n435), .Y(n334) );
  INV U706 ( .A(n636), .Y(n333) );
  MX2 U707 ( .A(n680), .B(\decider/posy_m_rex_top[1] ), .S0(n434), .Y(n636) );
  INV U708 ( .A(addrD[1]), .Y(n680) );
  INV U709 ( .A(n637), .Y(n332) );
  MX2 U710 ( .A(addrD[2]), .B(\decider/posy_m_rex_top[2] ), .S0(n435), .Y(n637) );
  INV U711 ( .A(n638), .Y(n331) );
  MX2 U712 ( .A(\decider/posy_m_obstacle_top [3]), .B(
        \decider/posy_m_rex_top[3] ), .S0(n434), .Y(n638) );
  INV U713 ( .A(n639), .Y(n330) );
  MX2 U714 ( .A(\decider/posy_m_obstacle_top [4]), .B(
        \decider/posy_m_rex_top[4] ), .S0(n435), .Y(n639) );
  INV U715 ( .A(n640), .Y(n329) );
  MX2 U716 ( .A(\decider/posy_m_obstacle_top [5]), .B(
        \decider/posy_m_rex_top[5] ), .S0(n434), .Y(n640) );
  NOR2B U717 ( .AN(rstn), .B(en_o), .Y(\driver/N96 ) );
  NOR2B U718 ( .AN(n435), .B(addrD[6]), .Y(\decider/N55 ) );
  NOR2B U719 ( .AN(addrD[10]), .B(n444), .Y(cs_o[3]) );
  NOR2B U720 ( .AN(addrD[10]), .B(addrD[9]), .Y(cs_o[2]) );
  NOR2B U721 ( .AN(n544), .B(n444), .Y(cs_o[1]) );
  NOR2B U722 ( .AN(\clock_divider/N17 ), .B(n433), .Y(\clock_divider/N30 ) );
  NOR2B U723 ( .AN(\clock_divider/N16 ), .B(n433), .Y(\clock_divider/N29 ) );
  NOR2B U724 ( .AN(\clock_divider/N15 ), .B(n433), .Y(\clock_divider/N28 ) );
  NOR2B U725 ( .AN(\clock_divider/N14 ), .B(n433), .Y(\clock_divider/N27 ) );
  NOR2B U726 ( .AN(\clock_divider/N13 ), .B(n433), .Y(\clock_divider/N26 ) );
  NOR2B U727 ( .AN(\clock_divider/N12 ), .B(n433), .Y(\clock_divider/N25 ) );
  NOR2B U728 ( .AN(\clock_divider/N11 ), .B(n433), .Y(\clock_divider/N24 ) );
  NOR2B U729 ( .AN(\clock_divider/N10 ), .B(n433), .Y(\clock_divider/N23 ) );
  NOR2B U730 ( .AN(\clock_divider/N9 ), .B(n433), .Y(\clock_divider/N22 ) );
  NOR2B U731 ( .AN(\clock_divider/N8 ), .B(n433), .Y(\clock_divider/N21 ) );
  NOR2B U732 ( .AN(\clock_divider/N7 ), .B(n433), .Y(\clock_divider/N20 ) );
  NOR2B U733 ( .AN(\clock_divider/N6 ), .B(n433), .Y(\clock_divider/N19 ) );
  NOR2B U734 ( .AN(n641), .B(n642), .Y(n635) );
  NAND4 U735 ( .A(\clock_divider/cnt5k[8] ), .B(\clock_divider/cnt5k[7] ), .C(
        \clock_divider/cnt5k[9] ), .D(n643), .Y(n642) );
  AND3 U736 ( .A(\clock_divider/cnt5k[1] ), .B(\clock_divider/cnt5k[12] ), .C(
        \clock_divider/cnt5k[2] ), .Y(n643) );
  NOR4BB U737 ( .AN(n644), .BN(\clock_divider/cnt5k[0] ), .C(
        \clock_divider/cnt5k[11] ), .D(\clock_divider/cnt5k[10] ), .Y(n641) );
  NOR4 U738 ( .A(\clock_divider/cnt5k[6] ), .B(\clock_divider/cnt5k[5] ), .C(
        \clock_divider/cnt5k[4] ), .D(\clock_divider/cnt5k[3] ), .Y(n644) );
  INV U739 ( .A(\clock_divider/cnt5k[0] ), .Y(\clock_divider/N18 ) );
  NOR2B U740 ( .AN(n677), .B(n434), .Y(\r62/ab[7][2] ) );
  NOR4BB U741 ( .AN(\decider/sub_45/carry[5] ), .BN(cs_o[0]), .C(addrD[8]), 
        .D(\sub_1_root_decider/sub_49/carry[6] ), .Y(n456) );
  NOR2B U742 ( .AN(n544), .B(addrD[9]), .Y(cs_o[0]) );
  INV U743 ( .A(addrD[10]), .Y(n544) );
  INV U744 ( .A(\r187/carry[8] ), .Y(n677) );
endmodule

